magic
tech gf180mcuC
magscale 1 10
timestamp 1670057553
<< metal1 >>
rect 60498 132638 60510 132690
rect 60562 132687 60574 132690
rect 61506 132687 61518 132690
rect 60562 132641 61518 132687
rect 60562 132638 60574 132641
rect 61506 132638 61518 132641
rect 61570 132638 61582 132690
rect 102834 132638 102846 132690
rect 102898 132687 102910 132690
rect 103730 132687 103742 132690
rect 102898 132641 103742 132687
rect 102898 132638 102910 132641
rect 103730 132638 103742 132641
rect 103794 132638 103806 132690
rect 1344 132522 118608 132556
rect 1344 132470 4478 132522
rect 4530 132470 4582 132522
rect 4634 132470 4686 132522
rect 4738 132470 35198 132522
rect 35250 132470 35302 132522
rect 35354 132470 35406 132522
rect 35458 132470 65918 132522
rect 65970 132470 66022 132522
rect 66074 132470 66126 132522
rect 66178 132470 96638 132522
rect 96690 132470 96742 132522
rect 96794 132470 96846 132522
rect 96898 132470 118608 132522
rect 1344 132436 118608 132470
rect 59838 132242 59890 132254
rect 22082 132190 22094 132242
rect 22146 132190 22158 132242
rect 59838 132178 59890 132190
rect 21410 132078 21422 132130
rect 21474 132078 21486 132130
rect 60834 132078 60846 132130
rect 60898 132078 60910 132130
rect 1822 132018 1874 132030
rect 1822 131954 1874 131966
rect 2494 132018 2546 132030
rect 2494 131954 2546 131966
rect 10334 132018 10386 132030
rect 10334 131954 10386 131966
rect 11678 132018 11730 132030
rect 11678 131954 11730 131966
rect 13582 132018 13634 132030
rect 13582 131954 13634 131966
rect 23774 132018 23826 132030
rect 23774 131954 23826 131966
rect 26462 132018 26514 132030
rect 26462 131954 26514 131966
rect 27806 132018 27858 132030
rect 27806 131954 27858 131966
rect 29822 132018 29874 132030
rect 29822 131954 29874 131966
rect 31166 132018 31218 132030
rect 31166 131954 31218 131966
rect 36318 132018 36370 132030
rect 36318 131954 36370 131966
rect 37214 132018 37266 132030
rect 37214 131954 37266 131966
rect 39902 132018 39954 132030
rect 39902 131954 39954 131966
rect 45950 132018 46002 132030
rect 45950 131954 46002 131966
rect 51326 132018 51378 132030
rect 51326 131954 51378 131966
rect 53342 132018 53394 132030
rect 53342 131954 53394 131966
rect 54686 132018 54738 132030
rect 54686 131954 54738 131966
rect 58718 132018 58770 132030
rect 58718 131954 58770 131966
rect 61518 132018 61570 132030
rect 61518 131954 61570 131966
rect 63422 132018 63474 132030
rect 63422 131954 63474 131966
rect 64766 132018 64818 132030
rect 64766 131954 64818 131966
rect 66110 132018 66162 132030
rect 66110 131954 66162 131966
rect 67454 132018 67506 132030
rect 67454 131954 67506 131966
rect 69470 132018 69522 132030
rect 69470 131954 69522 131966
rect 72382 132018 72434 132030
rect 72382 131954 72434 131966
rect 73502 132018 73554 132030
rect 73502 131954 73554 131966
rect 74846 132018 74898 132030
rect 74846 131954 74898 131966
rect 76302 132018 76354 132030
rect 76302 131954 76354 131966
rect 80894 132018 80946 132030
rect 80894 131954 80946 131966
rect 82238 132018 82290 132030
rect 82238 131954 82290 131966
rect 84254 132018 84306 132030
rect 84254 131954 84306 131966
rect 85598 132018 85650 132030
rect 85598 131954 85650 131966
rect 88286 132018 88338 132030
rect 88286 131954 88338 131966
rect 89630 132018 89682 132030
rect 89630 131954 89682 131966
rect 95902 132018 95954 132030
rect 95902 131954 95954 131966
rect 103742 132018 103794 132030
rect 103742 131954 103794 131966
rect 104414 132018 104466 132030
rect 104414 131954 104466 131966
rect 109118 132018 109170 132030
rect 109118 131954 109170 131966
rect 115502 132018 115554 132030
rect 115502 131954 115554 131966
rect 116510 132018 116562 132030
rect 116510 131954 116562 131966
rect 117294 132018 117346 132030
rect 117294 131954 117346 131966
rect 117854 132018 117906 132030
rect 117854 131954 117906 131966
rect 20638 131906 20690 131918
rect 20638 131842 20690 131854
rect 60622 131906 60674 131918
rect 60622 131842 60674 131854
rect 1344 131738 118608 131772
rect 1344 131686 19838 131738
rect 19890 131686 19942 131738
rect 19994 131686 20046 131738
rect 20098 131686 50558 131738
rect 50610 131686 50662 131738
rect 50714 131686 50766 131738
rect 50818 131686 81278 131738
rect 81330 131686 81382 131738
rect 81434 131686 81486 131738
rect 81538 131686 111998 131738
rect 112050 131686 112102 131738
rect 112154 131686 112206 131738
rect 112258 131686 118608 131738
rect 1344 131652 118608 131686
rect 1344 130954 118608 130988
rect 1344 130902 4478 130954
rect 4530 130902 4582 130954
rect 4634 130902 4686 130954
rect 4738 130902 35198 130954
rect 35250 130902 35302 130954
rect 35354 130902 35406 130954
rect 35458 130902 65918 130954
rect 65970 130902 66022 130954
rect 66074 130902 66126 130954
rect 66178 130902 96638 130954
rect 96690 130902 96742 130954
rect 96794 130902 96846 130954
rect 96898 130902 118608 130954
rect 1344 130868 118608 130902
rect 1822 130450 1874 130462
rect 1822 130386 1874 130398
rect 1344 130170 118608 130204
rect 1344 130118 19838 130170
rect 19890 130118 19942 130170
rect 19994 130118 20046 130170
rect 20098 130118 50558 130170
rect 50610 130118 50662 130170
rect 50714 130118 50766 130170
rect 50818 130118 81278 130170
rect 81330 130118 81382 130170
rect 81434 130118 81486 130170
rect 81538 130118 111998 130170
rect 112050 130118 112102 130170
rect 112154 130118 112206 130170
rect 112258 130118 118608 130170
rect 1344 130084 118608 130118
rect 1344 129386 118608 129420
rect 1344 129334 4478 129386
rect 4530 129334 4582 129386
rect 4634 129334 4686 129386
rect 4738 129334 35198 129386
rect 35250 129334 35302 129386
rect 35354 129334 35406 129386
rect 35458 129334 65918 129386
rect 65970 129334 66022 129386
rect 66074 129334 66126 129386
rect 66178 129334 96638 129386
rect 96690 129334 96742 129386
rect 96794 129334 96846 129386
rect 96898 129334 118608 129386
rect 1344 129300 118608 129334
rect 1344 128602 118608 128636
rect 1344 128550 19838 128602
rect 19890 128550 19942 128602
rect 19994 128550 20046 128602
rect 20098 128550 50558 128602
rect 50610 128550 50662 128602
rect 50714 128550 50766 128602
rect 50818 128550 81278 128602
rect 81330 128550 81382 128602
rect 81434 128550 81486 128602
rect 81538 128550 111998 128602
rect 112050 128550 112102 128602
rect 112154 128550 112206 128602
rect 112258 128550 118608 128602
rect 1344 128516 118608 128550
rect 1822 128322 1874 128334
rect 1822 128258 1874 128270
rect 1344 127818 118608 127852
rect 1344 127766 4478 127818
rect 4530 127766 4582 127818
rect 4634 127766 4686 127818
rect 4738 127766 35198 127818
rect 35250 127766 35302 127818
rect 35354 127766 35406 127818
rect 35458 127766 65918 127818
rect 65970 127766 66022 127818
rect 66074 127766 66126 127818
rect 66178 127766 96638 127818
rect 96690 127766 96742 127818
rect 96794 127766 96846 127818
rect 96898 127766 118608 127818
rect 1344 127732 118608 127766
rect 1822 127202 1874 127214
rect 1822 127138 1874 127150
rect 1344 127034 118608 127068
rect 1344 126982 19838 127034
rect 19890 126982 19942 127034
rect 19994 126982 20046 127034
rect 20098 126982 50558 127034
rect 50610 126982 50662 127034
rect 50714 126982 50766 127034
rect 50818 126982 81278 127034
rect 81330 126982 81382 127034
rect 81434 126982 81486 127034
rect 81538 126982 111998 127034
rect 112050 126982 112102 127034
rect 112154 126982 112206 127034
rect 112258 126982 118608 127034
rect 1344 126948 118608 126982
rect 118078 126754 118130 126766
rect 118078 126690 118130 126702
rect 1344 126250 118608 126284
rect 1344 126198 4478 126250
rect 4530 126198 4582 126250
rect 4634 126198 4686 126250
rect 4738 126198 35198 126250
rect 35250 126198 35302 126250
rect 35354 126198 35406 126250
rect 35458 126198 65918 126250
rect 65970 126198 66022 126250
rect 66074 126198 66126 126250
rect 66178 126198 96638 126250
rect 96690 126198 96742 126250
rect 96794 126198 96846 126250
rect 96898 126198 118608 126250
rect 1344 126164 118608 126198
rect 1344 125466 118608 125500
rect 1344 125414 19838 125466
rect 19890 125414 19942 125466
rect 19994 125414 20046 125466
rect 20098 125414 50558 125466
rect 50610 125414 50662 125466
rect 50714 125414 50766 125466
rect 50818 125414 81278 125466
rect 81330 125414 81382 125466
rect 81434 125414 81486 125466
rect 81538 125414 111998 125466
rect 112050 125414 112102 125466
rect 112154 125414 112206 125466
rect 112258 125414 118608 125466
rect 1344 125380 118608 125414
rect 1822 125186 1874 125198
rect 1822 125122 1874 125134
rect 1344 124682 118608 124716
rect 1344 124630 4478 124682
rect 4530 124630 4582 124682
rect 4634 124630 4686 124682
rect 4738 124630 35198 124682
rect 35250 124630 35302 124682
rect 35354 124630 35406 124682
rect 35458 124630 65918 124682
rect 65970 124630 66022 124682
rect 66074 124630 66126 124682
rect 66178 124630 96638 124682
rect 96690 124630 96742 124682
rect 96794 124630 96846 124682
rect 96898 124630 118608 124682
rect 1344 124596 118608 124630
rect 118078 124066 118130 124078
rect 118078 124002 118130 124014
rect 1344 123898 118608 123932
rect 1344 123846 19838 123898
rect 19890 123846 19942 123898
rect 19994 123846 20046 123898
rect 20098 123846 50558 123898
rect 50610 123846 50662 123898
rect 50714 123846 50766 123898
rect 50818 123846 81278 123898
rect 81330 123846 81382 123898
rect 81434 123846 81486 123898
rect 81538 123846 111998 123898
rect 112050 123846 112102 123898
rect 112154 123846 112206 123898
rect 112258 123846 118608 123898
rect 1344 123812 118608 123846
rect 1822 123618 1874 123630
rect 1822 123554 1874 123566
rect 1344 123114 118608 123148
rect 1344 123062 4478 123114
rect 4530 123062 4582 123114
rect 4634 123062 4686 123114
rect 4738 123062 35198 123114
rect 35250 123062 35302 123114
rect 35354 123062 35406 123114
rect 35458 123062 65918 123114
rect 65970 123062 66022 123114
rect 66074 123062 66126 123114
rect 66178 123062 96638 123114
rect 96690 123062 96742 123114
rect 96794 123062 96846 123114
rect 96898 123062 118608 123114
rect 1344 123028 118608 123062
rect 1344 122330 118608 122364
rect 1344 122278 19838 122330
rect 19890 122278 19942 122330
rect 19994 122278 20046 122330
rect 20098 122278 50558 122330
rect 50610 122278 50662 122330
rect 50714 122278 50766 122330
rect 50818 122278 81278 122330
rect 81330 122278 81382 122330
rect 81434 122278 81486 122330
rect 81538 122278 111998 122330
rect 112050 122278 112102 122330
rect 112154 122278 112206 122330
rect 112258 122278 118608 122330
rect 1344 122244 118608 122278
rect 1822 122050 1874 122062
rect 1822 121986 1874 121998
rect 1344 121546 118608 121580
rect 1344 121494 4478 121546
rect 4530 121494 4582 121546
rect 4634 121494 4686 121546
rect 4738 121494 35198 121546
rect 35250 121494 35302 121546
rect 35354 121494 35406 121546
rect 35458 121494 65918 121546
rect 65970 121494 66022 121546
rect 66074 121494 66126 121546
rect 66178 121494 96638 121546
rect 96690 121494 96742 121546
rect 96794 121494 96846 121546
rect 96898 121494 118608 121546
rect 1344 121460 118608 121494
rect 1344 120762 118608 120796
rect 1344 120710 19838 120762
rect 19890 120710 19942 120762
rect 19994 120710 20046 120762
rect 20098 120710 50558 120762
rect 50610 120710 50662 120762
rect 50714 120710 50766 120762
rect 50818 120710 81278 120762
rect 81330 120710 81382 120762
rect 81434 120710 81486 120762
rect 81538 120710 111998 120762
rect 112050 120710 112102 120762
rect 112154 120710 112206 120762
rect 112258 120710 118608 120762
rect 1344 120676 118608 120710
rect 1344 119978 118608 120012
rect 1344 119926 4478 119978
rect 4530 119926 4582 119978
rect 4634 119926 4686 119978
rect 4738 119926 35198 119978
rect 35250 119926 35302 119978
rect 35354 119926 35406 119978
rect 35458 119926 65918 119978
rect 65970 119926 66022 119978
rect 66074 119926 66126 119978
rect 66178 119926 96638 119978
rect 96690 119926 96742 119978
rect 96794 119926 96846 119978
rect 96898 119926 118608 119978
rect 1344 119892 118608 119926
rect 1344 119194 118608 119228
rect 1344 119142 19838 119194
rect 19890 119142 19942 119194
rect 19994 119142 20046 119194
rect 20098 119142 50558 119194
rect 50610 119142 50662 119194
rect 50714 119142 50766 119194
rect 50818 119142 81278 119194
rect 81330 119142 81382 119194
rect 81434 119142 81486 119194
rect 81538 119142 111998 119194
rect 112050 119142 112102 119194
rect 112154 119142 112206 119194
rect 112258 119142 118608 119194
rect 1344 119108 118608 119142
rect 1344 118410 118608 118444
rect 1344 118358 4478 118410
rect 4530 118358 4582 118410
rect 4634 118358 4686 118410
rect 4738 118358 35198 118410
rect 35250 118358 35302 118410
rect 35354 118358 35406 118410
rect 35458 118358 65918 118410
rect 65970 118358 66022 118410
rect 66074 118358 66126 118410
rect 66178 118358 96638 118410
rect 96690 118358 96742 118410
rect 96794 118358 96846 118410
rect 96898 118358 118608 118410
rect 1344 118324 118608 118358
rect 1344 117626 118608 117660
rect 1344 117574 19838 117626
rect 19890 117574 19942 117626
rect 19994 117574 20046 117626
rect 20098 117574 50558 117626
rect 50610 117574 50662 117626
rect 50714 117574 50766 117626
rect 50818 117574 81278 117626
rect 81330 117574 81382 117626
rect 81434 117574 81486 117626
rect 81538 117574 111998 117626
rect 112050 117574 112102 117626
rect 112154 117574 112206 117626
rect 112258 117574 118608 117626
rect 1344 117540 118608 117574
rect 1822 117346 1874 117358
rect 1822 117282 1874 117294
rect 1344 116842 118608 116876
rect 1344 116790 4478 116842
rect 4530 116790 4582 116842
rect 4634 116790 4686 116842
rect 4738 116790 35198 116842
rect 35250 116790 35302 116842
rect 35354 116790 35406 116842
rect 35458 116790 65918 116842
rect 65970 116790 66022 116842
rect 66074 116790 66126 116842
rect 66178 116790 96638 116842
rect 96690 116790 96742 116842
rect 96794 116790 96846 116842
rect 96898 116790 118608 116842
rect 1344 116756 118608 116790
rect 118078 116338 118130 116350
rect 118078 116274 118130 116286
rect 1344 116058 118608 116092
rect 1344 116006 19838 116058
rect 19890 116006 19942 116058
rect 19994 116006 20046 116058
rect 20098 116006 50558 116058
rect 50610 116006 50662 116058
rect 50714 116006 50766 116058
rect 50818 116006 81278 116058
rect 81330 116006 81382 116058
rect 81434 116006 81486 116058
rect 81538 116006 111998 116058
rect 112050 116006 112102 116058
rect 112154 116006 112206 116058
rect 112258 116006 118608 116058
rect 1344 115972 118608 116006
rect 118078 115778 118130 115790
rect 118078 115714 118130 115726
rect 1344 115274 118608 115308
rect 1344 115222 4478 115274
rect 4530 115222 4582 115274
rect 4634 115222 4686 115274
rect 4738 115222 35198 115274
rect 35250 115222 35302 115274
rect 35354 115222 35406 115274
rect 35458 115222 65918 115274
rect 65970 115222 66022 115274
rect 66074 115222 66126 115274
rect 66178 115222 96638 115274
rect 96690 115222 96742 115274
rect 96794 115222 96846 115274
rect 96898 115222 118608 115274
rect 1344 115188 118608 115222
rect 1344 114490 118608 114524
rect 1344 114438 19838 114490
rect 19890 114438 19942 114490
rect 19994 114438 20046 114490
rect 20098 114438 50558 114490
rect 50610 114438 50662 114490
rect 50714 114438 50766 114490
rect 50818 114438 81278 114490
rect 81330 114438 81382 114490
rect 81434 114438 81486 114490
rect 81538 114438 111998 114490
rect 112050 114438 112102 114490
rect 112154 114438 112206 114490
rect 112258 114438 118608 114490
rect 1344 114404 118608 114438
rect 118078 114322 118130 114334
rect 118078 114258 118130 114270
rect 1344 113706 118608 113740
rect 1344 113654 4478 113706
rect 4530 113654 4582 113706
rect 4634 113654 4686 113706
rect 4738 113654 35198 113706
rect 35250 113654 35302 113706
rect 35354 113654 35406 113706
rect 35458 113654 65918 113706
rect 65970 113654 66022 113706
rect 66074 113654 66126 113706
rect 66178 113654 96638 113706
rect 96690 113654 96742 113706
rect 96794 113654 96846 113706
rect 96898 113654 118608 113706
rect 1344 113620 118608 113654
rect 1344 112922 118608 112956
rect 1344 112870 19838 112922
rect 19890 112870 19942 112922
rect 19994 112870 20046 112922
rect 20098 112870 50558 112922
rect 50610 112870 50662 112922
rect 50714 112870 50766 112922
rect 50818 112870 81278 112922
rect 81330 112870 81382 112922
rect 81434 112870 81486 112922
rect 81538 112870 111998 112922
rect 112050 112870 112102 112922
rect 112154 112870 112206 112922
rect 112258 112870 118608 112922
rect 1344 112836 118608 112870
rect 1344 112138 118608 112172
rect 1344 112086 4478 112138
rect 4530 112086 4582 112138
rect 4634 112086 4686 112138
rect 4738 112086 35198 112138
rect 35250 112086 35302 112138
rect 35354 112086 35406 112138
rect 35458 112086 65918 112138
rect 65970 112086 66022 112138
rect 66074 112086 66126 112138
rect 66178 112086 96638 112138
rect 96690 112086 96742 112138
rect 96794 112086 96846 112138
rect 96898 112086 118608 112138
rect 1344 112052 118608 112086
rect 118078 111634 118130 111646
rect 118078 111570 118130 111582
rect 1822 111522 1874 111534
rect 1822 111458 1874 111470
rect 1344 111354 118608 111388
rect 1344 111302 19838 111354
rect 19890 111302 19942 111354
rect 19994 111302 20046 111354
rect 20098 111302 50558 111354
rect 50610 111302 50662 111354
rect 50714 111302 50766 111354
rect 50818 111302 81278 111354
rect 81330 111302 81382 111354
rect 81434 111302 81486 111354
rect 81538 111302 111998 111354
rect 112050 111302 112102 111354
rect 112154 111302 112206 111354
rect 112258 111302 118608 111354
rect 1344 111268 118608 111302
rect 118078 111074 118130 111086
rect 118078 111010 118130 111022
rect 1344 110570 118608 110604
rect 1344 110518 4478 110570
rect 4530 110518 4582 110570
rect 4634 110518 4686 110570
rect 4738 110518 35198 110570
rect 35250 110518 35302 110570
rect 35354 110518 35406 110570
rect 35458 110518 65918 110570
rect 65970 110518 66022 110570
rect 66074 110518 66126 110570
rect 66178 110518 96638 110570
rect 96690 110518 96742 110570
rect 96794 110518 96846 110570
rect 96898 110518 118608 110570
rect 1344 110484 118608 110518
rect 1822 109954 1874 109966
rect 1822 109890 1874 109902
rect 1344 109786 118608 109820
rect 1344 109734 19838 109786
rect 19890 109734 19942 109786
rect 19994 109734 20046 109786
rect 20098 109734 50558 109786
rect 50610 109734 50662 109786
rect 50714 109734 50766 109786
rect 50818 109734 81278 109786
rect 81330 109734 81382 109786
rect 81434 109734 81486 109786
rect 81538 109734 111998 109786
rect 112050 109734 112102 109786
rect 112154 109734 112206 109786
rect 112258 109734 118608 109786
rect 1344 109700 118608 109734
rect 1344 109002 118608 109036
rect 1344 108950 4478 109002
rect 4530 108950 4582 109002
rect 4634 108950 4686 109002
rect 4738 108950 35198 109002
rect 35250 108950 35302 109002
rect 35354 108950 35406 109002
rect 35458 108950 65918 109002
rect 65970 108950 66022 109002
rect 66074 108950 66126 109002
rect 66178 108950 96638 109002
rect 96690 108950 96742 109002
rect 96794 108950 96846 109002
rect 96898 108950 118608 109002
rect 1344 108916 118608 108950
rect 1344 108218 118608 108252
rect 1344 108166 19838 108218
rect 19890 108166 19942 108218
rect 19994 108166 20046 108218
rect 20098 108166 50558 108218
rect 50610 108166 50662 108218
rect 50714 108166 50766 108218
rect 50818 108166 81278 108218
rect 81330 108166 81382 108218
rect 81434 108166 81486 108218
rect 81538 108166 111998 108218
rect 112050 108166 112102 108218
rect 112154 108166 112206 108218
rect 112258 108166 118608 108218
rect 1344 108132 118608 108166
rect 118078 107938 118130 107950
rect 118078 107874 118130 107886
rect 1344 107434 118608 107468
rect 1344 107382 4478 107434
rect 4530 107382 4582 107434
rect 4634 107382 4686 107434
rect 4738 107382 35198 107434
rect 35250 107382 35302 107434
rect 35354 107382 35406 107434
rect 35458 107382 65918 107434
rect 65970 107382 66022 107434
rect 66074 107382 66126 107434
rect 66178 107382 96638 107434
rect 96690 107382 96742 107434
rect 96794 107382 96846 107434
rect 96898 107382 118608 107434
rect 1344 107348 118608 107382
rect 118078 106818 118130 106830
rect 118078 106754 118130 106766
rect 1344 106650 118608 106684
rect 1344 106598 19838 106650
rect 19890 106598 19942 106650
rect 19994 106598 20046 106650
rect 20098 106598 50558 106650
rect 50610 106598 50662 106650
rect 50714 106598 50766 106650
rect 50818 106598 81278 106650
rect 81330 106598 81382 106650
rect 81434 106598 81486 106650
rect 81538 106598 111998 106650
rect 112050 106598 112102 106650
rect 112154 106598 112206 106650
rect 112258 106598 118608 106650
rect 1344 106564 118608 106598
rect 1344 105866 118608 105900
rect 1344 105814 4478 105866
rect 4530 105814 4582 105866
rect 4634 105814 4686 105866
rect 4738 105814 35198 105866
rect 35250 105814 35302 105866
rect 35354 105814 35406 105866
rect 35458 105814 65918 105866
rect 65970 105814 66022 105866
rect 66074 105814 66126 105866
rect 66178 105814 96638 105866
rect 96690 105814 96742 105866
rect 96794 105814 96846 105866
rect 96898 105814 118608 105866
rect 1344 105780 118608 105814
rect 1822 105250 1874 105262
rect 1822 105186 1874 105198
rect 1344 105082 118608 105116
rect 1344 105030 19838 105082
rect 19890 105030 19942 105082
rect 19994 105030 20046 105082
rect 20098 105030 50558 105082
rect 50610 105030 50662 105082
rect 50714 105030 50766 105082
rect 50818 105030 81278 105082
rect 81330 105030 81382 105082
rect 81434 105030 81486 105082
rect 81538 105030 111998 105082
rect 112050 105030 112102 105082
rect 112154 105030 112206 105082
rect 112258 105030 118608 105082
rect 1344 104996 118608 105030
rect 1344 104298 118608 104332
rect 1344 104246 4478 104298
rect 4530 104246 4582 104298
rect 4634 104246 4686 104298
rect 4738 104246 35198 104298
rect 35250 104246 35302 104298
rect 35354 104246 35406 104298
rect 35458 104246 65918 104298
rect 65970 104246 66022 104298
rect 66074 104246 66126 104298
rect 66178 104246 96638 104298
rect 96690 104246 96742 104298
rect 96794 104246 96846 104298
rect 96898 104246 118608 104298
rect 1344 104212 118608 104246
rect 1344 103514 118608 103548
rect 1344 103462 19838 103514
rect 19890 103462 19942 103514
rect 19994 103462 20046 103514
rect 20098 103462 50558 103514
rect 50610 103462 50662 103514
rect 50714 103462 50766 103514
rect 50818 103462 81278 103514
rect 81330 103462 81382 103514
rect 81434 103462 81486 103514
rect 81538 103462 111998 103514
rect 112050 103462 112102 103514
rect 112154 103462 112206 103514
rect 112258 103462 118608 103514
rect 1344 103428 118608 103462
rect 118078 103234 118130 103246
rect 118078 103170 118130 103182
rect 1344 102730 118608 102764
rect 1344 102678 4478 102730
rect 4530 102678 4582 102730
rect 4634 102678 4686 102730
rect 4738 102678 35198 102730
rect 35250 102678 35302 102730
rect 35354 102678 35406 102730
rect 35458 102678 65918 102730
rect 65970 102678 66022 102730
rect 66074 102678 66126 102730
rect 66178 102678 96638 102730
rect 96690 102678 96742 102730
rect 96794 102678 96846 102730
rect 96898 102678 118608 102730
rect 1344 102644 118608 102678
rect 1344 101946 118608 101980
rect 1344 101894 19838 101946
rect 19890 101894 19942 101946
rect 19994 101894 20046 101946
rect 20098 101894 50558 101946
rect 50610 101894 50662 101946
rect 50714 101894 50766 101946
rect 50818 101894 81278 101946
rect 81330 101894 81382 101946
rect 81434 101894 81486 101946
rect 81538 101894 111998 101946
rect 112050 101894 112102 101946
rect 112154 101894 112206 101946
rect 112258 101894 118608 101946
rect 1344 101860 118608 101894
rect 1822 101666 1874 101678
rect 1822 101602 1874 101614
rect 1344 101162 118608 101196
rect 1344 101110 4478 101162
rect 4530 101110 4582 101162
rect 4634 101110 4686 101162
rect 4738 101110 35198 101162
rect 35250 101110 35302 101162
rect 35354 101110 35406 101162
rect 35458 101110 65918 101162
rect 65970 101110 66022 101162
rect 66074 101110 66126 101162
rect 66178 101110 96638 101162
rect 96690 101110 96742 101162
rect 96794 101110 96846 101162
rect 96898 101110 118608 101162
rect 1344 101076 118608 101110
rect 1344 100378 118608 100412
rect 1344 100326 19838 100378
rect 19890 100326 19942 100378
rect 19994 100326 20046 100378
rect 20098 100326 50558 100378
rect 50610 100326 50662 100378
rect 50714 100326 50766 100378
rect 50818 100326 81278 100378
rect 81330 100326 81382 100378
rect 81434 100326 81486 100378
rect 81538 100326 111998 100378
rect 112050 100326 112102 100378
rect 112154 100326 112206 100378
rect 112258 100326 118608 100378
rect 1344 100292 118608 100326
rect 1344 99594 118608 99628
rect 1344 99542 4478 99594
rect 4530 99542 4582 99594
rect 4634 99542 4686 99594
rect 4738 99542 35198 99594
rect 35250 99542 35302 99594
rect 35354 99542 35406 99594
rect 35458 99542 65918 99594
rect 65970 99542 66022 99594
rect 66074 99542 66126 99594
rect 66178 99542 96638 99594
rect 96690 99542 96742 99594
rect 96794 99542 96846 99594
rect 96898 99542 118608 99594
rect 1344 99508 118608 99542
rect 1344 98810 118608 98844
rect 1344 98758 19838 98810
rect 19890 98758 19942 98810
rect 19994 98758 20046 98810
rect 20098 98758 50558 98810
rect 50610 98758 50662 98810
rect 50714 98758 50766 98810
rect 50818 98758 81278 98810
rect 81330 98758 81382 98810
rect 81434 98758 81486 98810
rect 81538 98758 111998 98810
rect 112050 98758 112102 98810
rect 112154 98758 112206 98810
rect 112258 98758 118608 98810
rect 1344 98724 118608 98758
rect 118078 98530 118130 98542
rect 118078 98466 118130 98478
rect 1344 98026 118608 98060
rect 1344 97974 4478 98026
rect 4530 97974 4582 98026
rect 4634 97974 4686 98026
rect 4738 97974 35198 98026
rect 35250 97974 35302 98026
rect 35354 97974 35406 98026
rect 35458 97974 65918 98026
rect 65970 97974 66022 98026
rect 66074 97974 66126 98026
rect 66178 97974 96638 98026
rect 96690 97974 96742 98026
rect 96794 97974 96846 98026
rect 96898 97974 118608 98026
rect 1344 97940 118608 97974
rect 118078 97410 118130 97422
rect 118078 97346 118130 97358
rect 1344 97242 118608 97276
rect 1344 97190 19838 97242
rect 19890 97190 19942 97242
rect 19994 97190 20046 97242
rect 20098 97190 50558 97242
rect 50610 97190 50662 97242
rect 50714 97190 50766 97242
rect 50818 97190 81278 97242
rect 81330 97190 81382 97242
rect 81434 97190 81486 97242
rect 81538 97190 111998 97242
rect 112050 97190 112102 97242
rect 112154 97190 112206 97242
rect 112258 97190 118608 97242
rect 1344 97156 118608 97190
rect 1822 96962 1874 96974
rect 1822 96898 1874 96910
rect 1344 96458 118608 96492
rect 1344 96406 4478 96458
rect 4530 96406 4582 96458
rect 4634 96406 4686 96458
rect 4738 96406 35198 96458
rect 35250 96406 35302 96458
rect 35354 96406 35406 96458
rect 35458 96406 65918 96458
rect 65970 96406 66022 96458
rect 66074 96406 66126 96458
rect 66178 96406 96638 96458
rect 96690 96406 96742 96458
rect 96794 96406 96846 96458
rect 96898 96406 118608 96458
rect 1344 96372 118608 96406
rect 118078 95842 118130 95854
rect 118078 95778 118130 95790
rect 1344 95674 118608 95708
rect 1344 95622 19838 95674
rect 19890 95622 19942 95674
rect 19994 95622 20046 95674
rect 20098 95622 50558 95674
rect 50610 95622 50662 95674
rect 50714 95622 50766 95674
rect 50818 95622 81278 95674
rect 81330 95622 81382 95674
rect 81434 95622 81486 95674
rect 81538 95622 111998 95674
rect 112050 95622 112102 95674
rect 112154 95622 112206 95674
rect 112258 95622 118608 95674
rect 1344 95588 118608 95622
rect 1822 95394 1874 95406
rect 1822 95330 1874 95342
rect 1344 94890 118608 94924
rect 1344 94838 4478 94890
rect 4530 94838 4582 94890
rect 4634 94838 4686 94890
rect 4738 94838 35198 94890
rect 35250 94838 35302 94890
rect 35354 94838 35406 94890
rect 35458 94838 65918 94890
rect 65970 94838 66022 94890
rect 66074 94838 66126 94890
rect 66178 94838 96638 94890
rect 96690 94838 96742 94890
rect 96794 94838 96846 94890
rect 96898 94838 118608 94890
rect 1344 94804 118608 94838
rect 1344 94106 118608 94140
rect 1344 94054 19838 94106
rect 19890 94054 19942 94106
rect 19994 94054 20046 94106
rect 20098 94054 50558 94106
rect 50610 94054 50662 94106
rect 50714 94054 50766 94106
rect 50818 94054 81278 94106
rect 81330 94054 81382 94106
rect 81434 94054 81486 94106
rect 81538 94054 111998 94106
rect 112050 94054 112102 94106
rect 112154 94054 112206 94106
rect 112258 94054 118608 94106
rect 1344 94020 118608 94054
rect 1344 93322 118608 93356
rect 1344 93270 4478 93322
rect 4530 93270 4582 93322
rect 4634 93270 4686 93322
rect 4738 93270 35198 93322
rect 35250 93270 35302 93322
rect 35354 93270 35406 93322
rect 35458 93270 65918 93322
rect 65970 93270 66022 93322
rect 66074 93270 66126 93322
rect 66178 93270 96638 93322
rect 96690 93270 96742 93322
rect 96794 93270 96846 93322
rect 96898 93270 118608 93322
rect 1344 93236 118608 93270
rect 1822 92706 1874 92718
rect 1822 92642 1874 92654
rect 1344 92538 118608 92572
rect 1344 92486 19838 92538
rect 19890 92486 19942 92538
rect 19994 92486 20046 92538
rect 20098 92486 50558 92538
rect 50610 92486 50662 92538
rect 50714 92486 50766 92538
rect 50818 92486 81278 92538
rect 81330 92486 81382 92538
rect 81434 92486 81486 92538
rect 81538 92486 111998 92538
rect 112050 92486 112102 92538
rect 112154 92486 112206 92538
rect 112258 92486 118608 92538
rect 1344 92452 118608 92486
rect 1344 91754 118608 91788
rect 1344 91702 4478 91754
rect 4530 91702 4582 91754
rect 4634 91702 4686 91754
rect 4738 91702 35198 91754
rect 35250 91702 35302 91754
rect 35354 91702 35406 91754
rect 35458 91702 65918 91754
rect 65970 91702 66022 91754
rect 66074 91702 66126 91754
rect 66178 91702 96638 91754
rect 96690 91702 96742 91754
rect 96794 91702 96846 91754
rect 96898 91702 118608 91754
rect 1344 91668 118608 91702
rect 1822 91138 1874 91150
rect 1822 91074 1874 91086
rect 118078 91138 118130 91150
rect 118078 91074 118130 91086
rect 1344 90970 118608 91004
rect 1344 90918 19838 90970
rect 19890 90918 19942 90970
rect 19994 90918 20046 90970
rect 20098 90918 50558 90970
rect 50610 90918 50662 90970
rect 50714 90918 50766 90970
rect 50818 90918 81278 90970
rect 81330 90918 81382 90970
rect 81434 90918 81486 90970
rect 81538 90918 111998 90970
rect 112050 90918 112102 90970
rect 112154 90918 112206 90970
rect 112258 90918 118608 90970
rect 1344 90884 118608 90918
rect 2158 90690 2210 90702
rect 2158 90626 2210 90638
rect 1822 90578 1874 90590
rect 1822 90514 1874 90526
rect 1344 90186 118608 90220
rect 1344 90134 4478 90186
rect 4530 90134 4582 90186
rect 4634 90134 4686 90186
rect 4738 90134 35198 90186
rect 35250 90134 35302 90186
rect 35354 90134 35406 90186
rect 35458 90134 65918 90186
rect 65970 90134 66022 90186
rect 66074 90134 66126 90186
rect 66178 90134 96638 90186
rect 96690 90134 96742 90186
rect 96794 90134 96846 90186
rect 96898 90134 118608 90186
rect 1344 90100 118608 90134
rect 1822 89906 1874 89918
rect 1822 89842 1874 89854
rect 1344 89402 118608 89436
rect 1344 89350 19838 89402
rect 19890 89350 19942 89402
rect 19994 89350 20046 89402
rect 20098 89350 50558 89402
rect 50610 89350 50662 89402
rect 50714 89350 50766 89402
rect 50818 89350 81278 89402
rect 81330 89350 81382 89402
rect 81434 89350 81486 89402
rect 81538 89350 111998 89402
rect 112050 89350 112102 89402
rect 112154 89350 112206 89402
rect 112258 89350 118608 89402
rect 1344 89316 118608 89350
rect 1344 88618 118608 88652
rect 1344 88566 4478 88618
rect 4530 88566 4582 88618
rect 4634 88566 4686 88618
rect 4738 88566 35198 88618
rect 35250 88566 35302 88618
rect 35354 88566 35406 88618
rect 35458 88566 65918 88618
rect 65970 88566 66022 88618
rect 66074 88566 66126 88618
rect 66178 88566 96638 88618
rect 96690 88566 96742 88618
rect 96794 88566 96846 88618
rect 96898 88566 118608 88618
rect 1344 88532 118608 88566
rect 118078 88114 118130 88126
rect 118078 88050 118130 88062
rect 1344 87834 118608 87868
rect 1344 87782 19838 87834
rect 19890 87782 19942 87834
rect 19994 87782 20046 87834
rect 20098 87782 50558 87834
rect 50610 87782 50662 87834
rect 50714 87782 50766 87834
rect 50818 87782 81278 87834
rect 81330 87782 81382 87834
rect 81434 87782 81486 87834
rect 81538 87782 111998 87834
rect 112050 87782 112102 87834
rect 112154 87782 112206 87834
rect 112258 87782 118608 87834
rect 1344 87748 118608 87782
rect 1344 87050 118608 87084
rect 1344 86998 4478 87050
rect 4530 86998 4582 87050
rect 4634 86998 4686 87050
rect 4738 86998 35198 87050
rect 35250 86998 35302 87050
rect 35354 86998 35406 87050
rect 35458 86998 65918 87050
rect 65970 86998 66022 87050
rect 66074 86998 66126 87050
rect 66178 86998 96638 87050
rect 96690 86998 96742 87050
rect 96794 86998 96846 87050
rect 96898 86998 118608 87050
rect 1344 86964 118608 86998
rect 1344 86266 118608 86300
rect 1344 86214 19838 86266
rect 19890 86214 19942 86266
rect 19994 86214 20046 86266
rect 20098 86214 50558 86266
rect 50610 86214 50662 86266
rect 50714 86214 50766 86266
rect 50818 86214 81278 86266
rect 81330 86214 81382 86266
rect 81434 86214 81486 86266
rect 81538 86214 111998 86266
rect 112050 86214 112102 86266
rect 112154 86214 112206 86266
rect 112258 86214 118608 86266
rect 1344 86180 118608 86214
rect 1344 85482 118608 85516
rect 1344 85430 4478 85482
rect 4530 85430 4582 85482
rect 4634 85430 4686 85482
rect 4738 85430 35198 85482
rect 35250 85430 35302 85482
rect 35354 85430 35406 85482
rect 35458 85430 65918 85482
rect 65970 85430 66022 85482
rect 66074 85430 66126 85482
rect 66178 85430 96638 85482
rect 96690 85430 96742 85482
rect 96794 85430 96846 85482
rect 96898 85430 118608 85482
rect 1344 85396 118608 85430
rect 2818 85038 2830 85090
rect 2882 85038 2894 85090
rect 2146 84926 2158 84978
rect 2210 84926 2222 84978
rect 3502 84866 3554 84878
rect 3502 84802 3554 84814
rect 1344 84698 118608 84732
rect 1344 84646 19838 84698
rect 19890 84646 19942 84698
rect 19994 84646 20046 84698
rect 20098 84646 50558 84698
rect 50610 84646 50662 84698
rect 50714 84646 50766 84698
rect 50818 84646 81278 84698
rect 81330 84646 81382 84698
rect 81434 84646 81486 84698
rect 81538 84646 111998 84698
rect 112050 84646 112102 84698
rect 112154 84646 112206 84698
rect 112258 84646 118608 84698
rect 1344 84612 118608 84646
rect 118078 84418 118130 84430
rect 118078 84354 118130 84366
rect 1344 83914 118608 83948
rect 1344 83862 4478 83914
rect 4530 83862 4582 83914
rect 4634 83862 4686 83914
rect 4738 83862 35198 83914
rect 35250 83862 35302 83914
rect 35354 83862 35406 83914
rect 35458 83862 65918 83914
rect 65970 83862 66022 83914
rect 66074 83862 66126 83914
rect 66178 83862 96638 83914
rect 96690 83862 96742 83914
rect 96794 83862 96846 83914
rect 96898 83862 118608 83914
rect 1344 83828 118608 83862
rect 2494 83410 2546 83422
rect 2494 83346 2546 83358
rect 1822 83298 1874 83310
rect 1822 83234 1874 83246
rect 1344 83130 118608 83164
rect 1344 83078 19838 83130
rect 19890 83078 19942 83130
rect 19994 83078 20046 83130
rect 20098 83078 50558 83130
rect 50610 83078 50662 83130
rect 50714 83078 50766 83130
rect 50818 83078 81278 83130
rect 81330 83078 81382 83130
rect 81434 83078 81486 83130
rect 81538 83078 111998 83130
rect 112050 83078 112102 83130
rect 112154 83078 112206 83130
rect 112258 83078 118608 83130
rect 1344 83044 118608 83078
rect 118078 82850 118130 82862
rect 118078 82786 118130 82798
rect 1344 82346 118608 82380
rect 1344 82294 4478 82346
rect 4530 82294 4582 82346
rect 4634 82294 4686 82346
rect 4738 82294 35198 82346
rect 35250 82294 35302 82346
rect 35354 82294 35406 82346
rect 35458 82294 65918 82346
rect 65970 82294 66022 82346
rect 66074 82294 66126 82346
rect 66178 82294 96638 82346
rect 96690 82294 96742 82346
rect 96794 82294 96846 82346
rect 96898 82294 118608 82346
rect 1344 82260 118608 82294
rect 1344 81562 118608 81596
rect 1344 81510 19838 81562
rect 19890 81510 19942 81562
rect 19994 81510 20046 81562
rect 20098 81510 50558 81562
rect 50610 81510 50662 81562
rect 50714 81510 50766 81562
rect 50818 81510 81278 81562
rect 81330 81510 81382 81562
rect 81434 81510 81486 81562
rect 81538 81510 111998 81562
rect 112050 81510 112102 81562
rect 112154 81510 112206 81562
rect 112258 81510 118608 81562
rect 1344 81476 118608 81510
rect 1344 80778 118608 80812
rect 1344 80726 4478 80778
rect 4530 80726 4582 80778
rect 4634 80726 4686 80778
rect 4738 80726 35198 80778
rect 35250 80726 35302 80778
rect 35354 80726 35406 80778
rect 35458 80726 65918 80778
rect 65970 80726 66022 80778
rect 66074 80726 66126 80778
rect 66178 80726 96638 80778
rect 96690 80726 96742 80778
rect 96794 80726 96846 80778
rect 96898 80726 118608 80778
rect 1344 80692 118608 80726
rect 1344 79994 118608 80028
rect 1344 79942 19838 79994
rect 19890 79942 19942 79994
rect 19994 79942 20046 79994
rect 20098 79942 50558 79994
rect 50610 79942 50662 79994
rect 50714 79942 50766 79994
rect 50818 79942 81278 79994
rect 81330 79942 81382 79994
rect 81434 79942 81486 79994
rect 81538 79942 111998 79994
rect 112050 79942 112102 79994
rect 112154 79942 112206 79994
rect 112258 79942 118608 79994
rect 1344 79908 118608 79942
rect 118078 79714 118130 79726
rect 118078 79650 118130 79662
rect 1344 79210 118608 79244
rect 1344 79158 4478 79210
rect 4530 79158 4582 79210
rect 4634 79158 4686 79210
rect 4738 79158 35198 79210
rect 35250 79158 35302 79210
rect 35354 79158 35406 79210
rect 35458 79158 65918 79210
rect 65970 79158 66022 79210
rect 66074 79158 66126 79210
rect 66178 79158 96638 79210
rect 96690 79158 96742 79210
rect 96794 79158 96846 79210
rect 96898 79158 118608 79210
rect 1344 79124 118608 79158
rect 1344 78426 118608 78460
rect 1344 78374 19838 78426
rect 19890 78374 19942 78426
rect 19994 78374 20046 78426
rect 20098 78374 50558 78426
rect 50610 78374 50662 78426
rect 50714 78374 50766 78426
rect 50818 78374 81278 78426
rect 81330 78374 81382 78426
rect 81434 78374 81486 78426
rect 81538 78374 111998 78426
rect 112050 78374 112102 78426
rect 112154 78374 112206 78426
rect 112258 78374 118608 78426
rect 1344 78340 118608 78374
rect 2158 78146 2210 78158
rect 2158 78082 2210 78094
rect 1822 78034 1874 78046
rect 1822 77970 1874 77982
rect 1344 77642 118608 77676
rect 1344 77590 4478 77642
rect 4530 77590 4582 77642
rect 4634 77590 4686 77642
rect 4738 77590 35198 77642
rect 35250 77590 35302 77642
rect 35354 77590 35406 77642
rect 35458 77590 65918 77642
rect 65970 77590 66022 77642
rect 66074 77590 66126 77642
rect 66178 77590 96638 77642
rect 96690 77590 96742 77642
rect 96794 77590 96846 77642
rect 96898 77590 118608 77642
rect 1344 77556 118608 77590
rect 1822 77362 1874 77374
rect 1822 77298 1874 77310
rect 118078 77026 118130 77038
rect 118078 76962 118130 76974
rect 1344 76858 118608 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 81278 76858
rect 81330 76806 81382 76858
rect 81434 76806 81486 76858
rect 81538 76806 111998 76858
rect 112050 76806 112102 76858
rect 112154 76806 112206 76858
rect 112258 76806 118608 76858
rect 1344 76772 118608 76806
rect 1344 76074 118608 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 96638 76074
rect 96690 76022 96742 76074
rect 96794 76022 96846 76074
rect 96898 76022 118608 76074
rect 1344 75988 118608 76022
rect 1344 75290 118608 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 81278 75290
rect 81330 75238 81382 75290
rect 81434 75238 81486 75290
rect 81538 75238 111998 75290
rect 112050 75238 112102 75290
rect 112154 75238 112206 75290
rect 112258 75238 118608 75290
rect 1344 75204 118608 75238
rect 1344 74506 118608 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 96638 74506
rect 96690 74454 96742 74506
rect 96794 74454 96846 74506
rect 96898 74454 118608 74506
rect 1344 74420 118608 74454
rect 118078 73890 118130 73902
rect 118078 73826 118130 73838
rect 1344 73722 118608 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 81278 73722
rect 81330 73670 81382 73722
rect 81434 73670 81486 73722
rect 81538 73670 111998 73722
rect 112050 73670 112102 73722
rect 112154 73670 112206 73722
rect 112258 73670 118608 73722
rect 1344 73636 118608 73670
rect 1822 73442 1874 73454
rect 1822 73378 1874 73390
rect 1344 72938 118608 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 96638 72938
rect 96690 72886 96742 72938
rect 96794 72886 96846 72938
rect 96898 72886 118608 72938
rect 1344 72852 118608 72886
rect 1344 72154 118608 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 81278 72154
rect 81330 72102 81382 72154
rect 81434 72102 81486 72154
rect 81538 72102 111998 72154
rect 112050 72102 112102 72154
rect 112154 72102 112206 72154
rect 112258 72102 118608 72154
rect 1344 72068 118608 72102
rect 1344 71370 118608 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 96638 71370
rect 96690 71318 96742 71370
rect 96794 71318 96846 71370
rect 96898 71318 118608 71370
rect 1344 71284 118608 71318
rect 1344 70586 118608 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 81278 70586
rect 81330 70534 81382 70586
rect 81434 70534 81486 70586
rect 81538 70534 111998 70586
rect 112050 70534 112102 70586
rect 112154 70534 112206 70586
rect 112258 70534 118608 70586
rect 1344 70500 118608 70534
rect 1344 69802 118608 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 96638 69802
rect 96690 69750 96742 69802
rect 96794 69750 96846 69802
rect 96898 69750 118608 69802
rect 1344 69716 118608 69750
rect 118078 69298 118130 69310
rect 118078 69234 118130 69246
rect 1344 69018 118608 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 81278 69018
rect 81330 68966 81382 69018
rect 81434 68966 81486 69018
rect 81538 68966 111998 69018
rect 112050 68966 112102 69018
rect 112154 68966 112206 69018
rect 112258 68966 118608 69018
rect 1344 68932 118608 68966
rect 3166 68850 3218 68862
rect 3166 68786 3218 68798
rect 20078 68850 20130 68862
rect 20078 68786 20130 68798
rect 2606 68738 2658 68750
rect 2606 68674 2658 68686
rect 118078 68738 118130 68750
rect 118078 68674 118130 68686
rect 19966 68514 20018 68526
rect 19966 68450 20018 68462
rect 20638 68514 20690 68526
rect 20638 68450 20690 68462
rect 2718 68402 2770 68414
rect 2718 68338 2770 68350
rect 1344 68234 118608 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 96638 68234
rect 96690 68182 96742 68234
rect 96794 68182 96846 68234
rect 96898 68182 118608 68234
rect 1344 68148 118608 68182
rect 60062 67954 60114 67966
rect 60062 67890 60114 67902
rect 3390 67842 3442 67854
rect 3390 67778 3442 67790
rect 4062 67842 4114 67854
rect 4062 67778 4114 67790
rect 59614 67842 59666 67854
rect 59614 67778 59666 67790
rect 2046 67730 2098 67742
rect 2046 67666 2098 67678
rect 2494 67730 2546 67742
rect 2494 67666 2546 67678
rect 2830 67730 2882 67742
rect 2830 67666 2882 67678
rect 3502 67618 3554 67630
rect 3502 67554 3554 67566
rect 3726 67618 3778 67630
rect 3726 67554 3778 67566
rect 59278 67618 59330 67630
rect 59278 67554 59330 67566
rect 118078 67618 118130 67630
rect 118078 67554 118130 67566
rect 1344 67450 118608 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 81278 67450
rect 81330 67398 81382 67450
rect 81434 67398 81486 67450
rect 81538 67398 111998 67450
rect 112050 67398 112102 67450
rect 112154 67398 112206 67450
rect 112258 67398 118608 67450
rect 1344 67364 118608 67398
rect 6302 67170 6354 67182
rect 6302 67106 6354 67118
rect 1922 67006 1934 67058
rect 1986 67006 1998 67058
rect 2258 67006 2270 67058
rect 2322 67006 2334 67058
rect 4610 67006 4622 67058
rect 4674 67006 4686 67058
rect 5058 67006 5070 67058
rect 5122 67006 5134 67058
rect 5854 66834 5906 66846
rect 5854 66770 5906 66782
rect 1344 66666 118608 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 96638 66666
rect 96690 66614 96742 66666
rect 96794 66614 96846 66666
rect 96898 66614 118608 66666
rect 1344 66580 118608 66614
rect 1822 66274 1874 66286
rect 1822 66210 1874 66222
rect 2158 66162 2210 66174
rect 2158 66098 2210 66110
rect 1344 65882 118608 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 81278 65882
rect 81330 65830 81382 65882
rect 81434 65830 81486 65882
rect 81538 65830 111998 65882
rect 112050 65830 112102 65882
rect 112154 65830 112206 65882
rect 112258 65830 118608 65882
rect 1344 65796 118608 65830
rect 1822 65714 1874 65726
rect 1822 65650 1874 65662
rect 1344 65098 118608 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 96638 65098
rect 96690 65046 96742 65098
rect 96794 65046 96846 65098
rect 96898 65046 118608 65098
rect 1344 65012 118608 65046
rect 1822 64482 1874 64494
rect 1822 64418 1874 64430
rect 1344 64314 118608 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 81278 64314
rect 81330 64262 81382 64314
rect 81434 64262 81486 64314
rect 81538 64262 111998 64314
rect 112050 64262 112102 64314
rect 112154 64262 112206 64314
rect 112258 64262 118608 64314
rect 1344 64228 118608 64262
rect 1344 63530 118608 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 96638 63530
rect 96690 63478 96742 63530
rect 96794 63478 96846 63530
rect 96898 63478 118608 63530
rect 1344 63444 118608 63478
rect 1344 62746 118608 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 81278 62746
rect 81330 62694 81382 62746
rect 81434 62694 81486 62746
rect 81538 62694 111998 62746
rect 112050 62694 112102 62746
rect 112154 62694 112206 62746
rect 112258 62694 118608 62746
rect 1344 62660 118608 62694
rect 1344 61962 118608 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 96638 61962
rect 96690 61910 96742 61962
rect 96794 61910 96846 61962
rect 96898 61910 118608 61962
rect 1344 61876 118608 61910
rect 1822 61346 1874 61358
rect 1822 61282 1874 61294
rect 1344 61178 118608 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 81278 61178
rect 81330 61126 81382 61178
rect 81434 61126 81486 61178
rect 81538 61126 111998 61178
rect 112050 61126 112102 61178
rect 112154 61126 112206 61178
rect 112258 61126 118608 61178
rect 1344 61092 118608 61126
rect 118078 60898 118130 60910
rect 118078 60834 118130 60846
rect 1344 60394 118608 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 96638 60394
rect 96690 60342 96742 60394
rect 96794 60342 96846 60394
rect 96898 60342 118608 60394
rect 1344 60308 118608 60342
rect 118078 59890 118130 59902
rect 118078 59826 118130 59838
rect 1344 59610 118608 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 81278 59610
rect 81330 59558 81382 59610
rect 81434 59558 81486 59610
rect 81538 59558 111998 59610
rect 112050 59558 112102 59610
rect 112154 59558 112206 59610
rect 112258 59558 118608 59610
rect 1344 59524 118608 59558
rect 118078 59330 118130 59342
rect 118078 59266 118130 59278
rect 1344 58826 118608 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 96638 58826
rect 96690 58774 96742 58826
rect 96794 58774 96846 58826
rect 96898 58774 118608 58826
rect 1344 58740 118608 58774
rect 1822 58210 1874 58222
rect 1822 58146 1874 58158
rect 1344 58042 118608 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 81278 58042
rect 81330 57990 81382 58042
rect 81434 57990 81486 58042
rect 81538 57990 111998 58042
rect 112050 57990 112102 58042
rect 112154 57990 112206 58042
rect 112258 57990 118608 58042
rect 1344 57956 118608 57990
rect 118078 57762 118130 57774
rect 118078 57698 118130 57710
rect 1344 57258 118608 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 96638 57258
rect 96690 57206 96742 57258
rect 96794 57206 96846 57258
rect 96898 57206 118608 57258
rect 1344 57172 118608 57206
rect 1344 56474 118608 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 81278 56474
rect 81330 56422 81382 56474
rect 81434 56422 81486 56474
rect 81538 56422 111998 56474
rect 112050 56422 112102 56474
rect 112154 56422 112206 56474
rect 112258 56422 118608 56474
rect 1344 56388 118608 56422
rect 1344 55690 118608 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 96638 55690
rect 96690 55638 96742 55690
rect 96794 55638 96846 55690
rect 96898 55638 118608 55690
rect 1344 55604 118608 55638
rect 1344 54906 118608 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 81278 54906
rect 81330 54854 81382 54906
rect 81434 54854 81486 54906
rect 81538 54854 111998 54906
rect 112050 54854 112102 54906
rect 112154 54854 112206 54906
rect 112258 54854 118608 54906
rect 1344 54820 118608 54854
rect 1344 54122 118608 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 96638 54122
rect 96690 54070 96742 54122
rect 96794 54070 96846 54122
rect 96898 54070 118608 54122
rect 1344 54036 118608 54070
rect 118078 53506 118130 53518
rect 118078 53442 118130 53454
rect 1344 53338 118608 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 81278 53338
rect 81330 53286 81382 53338
rect 81434 53286 81486 53338
rect 81538 53286 111998 53338
rect 112050 53286 112102 53338
rect 112154 53286 112206 53338
rect 112258 53286 118608 53338
rect 1344 53252 118608 53286
rect 2158 53170 2210 53182
rect 2158 53106 2210 53118
rect 118078 53058 118130 53070
rect 118078 52994 118130 53006
rect 1822 52946 1874 52958
rect 1822 52882 1874 52894
rect 1344 52554 118608 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 96638 52554
rect 96690 52502 96742 52554
rect 96794 52502 96846 52554
rect 96898 52502 118608 52554
rect 1344 52468 118608 52502
rect 1822 52274 1874 52286
rect 1822 52210 1874 52222
rect 1344 51770 118608 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 81278 51770
rect 81330 51718 81382 51770
rect 81434 51718 81486 51770
rect 81538 51718 111998 51770
rect 112050 51718 112102 51770
rect 112154 51718 112206 51770
rect 112258 51718 118608 51770
rect 1344 51684 118608 51718
rect 1344 50986 118608 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 96638 50986
rect 96690 50934 96742 50986
rect 96794 50934 96846 50986
rect 96898 50934 118608 50986
rect 1344 50900 118608 50934
rect 1344 50202 118608 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 81278 50202
rect 81330 50150 81382 50202
rect 81434 50150 81486 50202
rect 81538 50150 111998 50202
rect 112050 50150 112102 50202
rect 112154 50150 112206 50202
rect 112258 50150 118608 50202
rect 1344 50116 118608 50150
rect 1822 49922 1874 49934
rect 1822 49858 1874 49870
rect 1344 49418 118608 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 96638 49418
rect 96690 49366 96742 49418
rect 96794 49366 96846 49418
rect 96898 49366 118608 49418
rect 1344 49332 118608 49366
rect 1344 48634 118608 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 81278 48634
rect 81330 48582 81382 48634
rect 81434 48582 81486 48634
rect 81538 48582 111998 48634
rect 112050 48582 112102 48634
rect 112154 48582 112206 48634
rect 112258 48582 118608 48634
rect 1344 48548 118608 48582
rect 3042 48190 3054 48242
rect 3106 48190 3118 48242
rect 3502 48130 3554 48142
rect 2034 48078 2046 48130
rect 2098 48078 2110 48130
rect 3502 48066 3554 48078
rect 1344 47850 118608 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 96638 47850
rect 96690 47798 96742 47850
rect 96794 47798 96846 47850
rect 96898 47798 118608 47850
rect 1344 47764 118608 47798
rect 118078 47234 118130 47246
rect 118078 47170 118130 47182
rect 1344 47066 118608 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 81278 47066
rect 81330 47014 81382 47066
rect 81434 47014 81486 47066
rect 81538 47014 111998 47066
rect 112050 47014 112102 47066
rect 112154 47014 112206 47066
rect 112258 47014 118608 47066
rect 1344 46980 118608 47014
rect 1822 46786 1874 46798
rect 1822 46722 1874 46734
rect 1344 46282 118608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 96638 46282
rect 96690 46230 96742 46282
rect 96794 46230 96846 46282
rect 96898 46230 118608 46282
rect 1344 46196 118608 46230
rect 1922 45838 1934 45890
rect 1986 45838 1998 45890
rect 2158 45666 2210 45678
rect 2158 45602 2210 45614
rect 2606 45666 2658 45678
rect 2606 45602 2658 45614
rect 118078 45666 118130 45678
rect 118078 45602 118130 45614
rect 1344 45498 118608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 81278 45498
rect 81330 45446 81382 45498
rect 81434 45446 81486 45498
rect 81538 45446 111998 45498
rect 112050 45446 112102 45498
rect 112154 45446 112206 45498
rect 112258 45446 118608 45498
rect 1344 45412 118608 45446
rect 2158 45330 2210 45342
rect 2158 45266 2210 45278
rect 1822 45106 1874 45118
rect 1822 45042 1874 45054
rect 1344 44714 118608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 96638 44714
rect 96690 44662 96742 44714
rect 96794 44662 96846 44714
rect 96898 44662 118608 44714
rect 1344 44628 118608 44662
rect 1822 44434 1874 44446
rect 1822 44370 1874 44382
rect 118078 44098 118130 44110
rect 118078 44034 118130 44046
rect 1344 43930 118608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 81278 43930
rect 81330 43878 81382 43930
rect 81434 43878 81486 43930
rect 81538 43878 111998 43930
rect 112050 43878 112102 43930
rect 112154 43878 112206 43930
rect 112258 43878 118608 43930
rect 1344 43844 118608 43878
rect 1344 43146 118608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 96638 43146
rect 96690 43094 96742 43146
rect 96794 43094 96846 43146
rect 96898 43094 118608 43146
rect 1344 43060 118608 43094
rect 1344 42362 118608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 81278 42362
rect 81330 42310 81382 42362
rect 81434 42310 81486 42362
rect 81538 42310 111998 42362
rect 112050 42310 112102 42362
rect 112154 42310 112206 42362
rect 112258 42310 118608 42362
rect 1344 42276 118608 42310
rect 1822 42082 1874 42094
rect 1822 42018 1874 42030
rect 1344 41578 118608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 96638 41578
rect 96690 41526 96742 41578
rect 96794 41526 96846 41578
rect 96898 41526 118608 41578
rect 1344 41492 118608 41526
rect 59950 41074 60002 41086
rect 59950 41010 60002 41022
rect 118078 41074 118130 41086
rect 118078 41010 118130 41022
rect 1822 40962 1874 40974
rect 1822 40898 1874 40910
rect 59390 40962 59442 40974
rect 59390 40898 59442 40910
rect 60286 40962 60338 40974
rect 60286 40898 60338 40910
rect 1344 40794 118608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 81278 40794
rect 81330 40742 81382 40794
rect 81434 40742 81486 40794
rect 81538 40742 111998 40794
rect 112050 40742 112102 40794
rect 112154 40742 112206 40794
rect 112258 40742 118608 40794
rect 1344 40708 118608 40742
rect 1344 40010 118608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 96638 40010
rect 96690 39958 96742 40010
rect 96794 39958 96846 40010
rect 96898 39958 118608 40010
rect 1344 39924 118608 39958
rect 1822 39394 1874 39406
rect 1822 39330 1874 39342
rect 1344 39226 118608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 81278 39226
rect 81330 39174 81382 39226
rect 81434 39174 81486 39226
rect 81538 39174 111998 39226
rect 112050 39174 112102 39226
rect 112154 39174 112206 39226
rect 112258 39174 118608 39226
rect 1344 39140 118608 39174
rect 118078 38946 118130 38958
rect 118078 38882 118130 38894
rect 1344 38442 118608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 96638 38442
rect 96690 38390 96742 38442
rect 96794 38390 96846 38442
rect 96898 38390 118608 38442
rect 1344 38356 118608 38390
rect 1344 37658 118608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 81278 37658
rect 81330 37606 81382 37658
rect 81434 37606 81486 37658
rect 81538 37606 111998 37658
rect 112050 37606 112102 37658
rect 112154 37606 112206 37658
rect 112258 37606 118608 37658
rect 1344 37572 118608 37606
rect 1822 37378 1874 37390
rect 1822 37314 1874 37326
rect 1344 36874 118608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 96638 36874
rect 96690 36822 96742 36874
rect 96794 36822 96846 36874
rect 96898 36822 118608 36874
rect 1344 36788 118608 36822
rect 1822 36258 1874 36270
rect 1822 36194 1874 36206
rect 1344 36090 118608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 81278 36090
rect 81330 36038 81382 36090
rect 81434 36038 81486 36090
rect 81538 36038 111998 36090
rect 112050 36038 112102 36090
rect 112154 36038 112206 36090
rect 112258 36038 118608 36090
rect 1344 36004 118608 36038
rect 117730 35758 117742 35810
rect 117794 35758 117806 35810
rect 116834 35646 116846 35698
rect 116898 35646 116910 35698
rect 116286 35586 116338 35598
rect 116286 35522 116338 35534
rect 1344 35306 118608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 96638 35306
rect 96690 35254 96742 35306
rect 96794 35254 96846 35306
rect 96898 35254 118608 35306
rect 1344 35220 118608 35254
rect 1344 34522 118608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 81278 34522
rect 81330 34470 81382 34522
rect 81434 34470 81486 34522
rect 81538 34470 111998 34522
rect 112050 34470 112102 34522
rect 112154 34470 112206 34522
rect 112258 34470 118608 34522
rect 1344 34436 118608 34470
rect 1344 33738 118608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 96638 33738
rect 96690 33686 96742 33738
rect 96794 33686 96846 33738
rect 96898 33686 118608 33738
rect 1344 33652 118608 33686
rect 1822 33122 1874 33134
rect 1822 33058 1874 33070
rect 1344 32954 118608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 81278 32954
rect 81330 32902 81382 32954
rect 81434 32902 81486 32954
rect 81538 32902 111998 32954
rect 112050 32902 112102 32954
rect 112154 32902 112206 32954
rect 112258 32902 118608 32954
rect 1344 32868 118608 32902
rect 1344 32170 118608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 96638 32170
rect 96690 32118 96742 32170
rect 96794 32118 96846 32170
rect 96898 32118 118608 32170
rect 1344 32084 118608 32118
rect 118078 31554 118130 31566
rect 118078 31490 118130 31502
rect 1344 31386 118608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 81278 31386
rect 81330 31334 81382 31386
rect 81434 31334 81486 31386
rect 81538 31334 111998 31386
rect 112050 31334 112102 31386
rect 112154 31334 112206 31386
rect 112258 31334 118608 31386
rect 1344 31300 118608 31334
rect 1344 30602 118608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 96638 30602
rect 96690 30550 96742 30602
rect 96794 30550 96846 30602
rect 96898 30550 118608 30602
rect 1344 30516 118608 30550
rect 1822 29986 1874 29998
rect 1822 29922 1874 29934
rect 1344 29818 118608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 81278 29818
rect 81330 29766 81382 29818
rect 81434 29766 81486 29818
rect 81538 29766 111998 29818
rect 112050 29766 112102 29818
rect 112154 29766 112206 29818
rect 112258 29766 118608 29818
rect 1344 29732 118608 29766
rect 118078 29538 118130 29550
rect 118078 29474 118130 29486
rect 1344 29034 118608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 96638 29034
rect 96690 28982 96742 29034
rect 96794 28982 96846 29034
rect 96898 28982 118608 29034
rect 1344 28948 118608 28982
rect 1344 28250 118608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 81278 28250
rect 81330 28198 81382 28250
rect 81434 28198 81486 28250
rect 81538 28198 111998 28250
rect 112050 28198 112102 28250
rect 112154 28198 112206 28250
rect 112258 28198 118608 28250
rect 1344 28164 118608 28198
rect 1344 27466 118608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 96638 27466
rect 96690 27414 96742 27466
rect 96794 27414 96846 27466
rect 96898 27414 118608 27466
rect 1344 27380 118608 27414
rect 118078 26850 118130 26862
rect 118078 26786 118130 26798
rect 1344 26682 118608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 81278 26682
rect 81330 26630 81382 26682
rect 81434 26630 81486 26682
rect 81538 26630 111998 26682
rect 112050 26630 112102 26682
rect 112154 26630 112206 26682
rect 112258 26630 118608 26682
rect 1344 26596 118608 26630
rect 1822 26402 1874 26414
rect 1822 26338 1874 26350
rect 1344 25898 118608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 96638 25898
rect 96690 25846 96742 25898
rect 96794 25846 96846 25898
rect 96898 25846 118608 25898
rect 1344 25812 118608 25846
rect 118078 25282 118130 25294
rect 118078 25218 118130 25230
rect 1344 25114 118608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 81278 25114
rect 81330 25062 81382 25114
rect 81434 25062 81486 25114
rect 81538 25062 111998 25114
rect 112050 25062 112102 25114
rect 112154 25062 112206 25114
rect 112258 25062 118608 25114
rect 1344 25028 118608 25062
rect 1344 24330 118608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 96638 24330
rect 96690 24278 96742 24330
rect 96794 24278 96846 24330
rect 96898 24278 118608 24330
rect 1344 24244 118608 24278
rect 1344 23546 118608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 81278 23546
rect 81330 23494 81382 23546
rect 81434 23494 81486 23546
rect 81538 23494 111998 23546
rect 112050 23494 112102 23546
rect 112154 23494 112206 23546
rect 112258 23494 118608 23546
rect 1344 23460 118608 23494
rect 1822 23266 1874 23278
rect 1822 23202 1874 23214
rect 118078 23266 118130 23278
rect 118078 23202 118130 23214
rect 1344 22762 118608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 96638 22762
rect 96690 22710 96742 22762
rect 96794 22710 96846 22762
rect 96898 22710 118608 22762
rect 1344 22676 118608 22710
rect 1344 21978 118608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 81278 21978
rect 81330 21926 81382 21978
rect 81434 21926 81486 21978
rect 81538 21926 111998 21978
rect 112050 21926 112102 21978
rect 112154 21926 112206 21978
rect 112258 21926 118608 21978
rect 1344 21892 118608 21926
rect 1822 21698 1874 21710
rect 1822 21634 1874 21646
rect 1344 21194 118608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 96638 21194
rect 96690 21142 96742 21194
rect 96794 21142 96846 21194
rect 96898 21142 118608 21194
rect 1344 21108 118608 21142
rect 118078 20578 118130 20590
rect 118078 20514 118130 20526
rect 1344 20410 118608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 81278 20410
rect 81330 20358 81382 20410
rect 81434 20358 81486 20410
rect 81538 20358 111998 20410
rect 112050 20358 112102 20410
rect 112154 20358 112206 20410
rect 112258 20358 118608 20410
rect 1344 20324 118608 20358
rect 1344 19626 118608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 96638 19626
rect 96690 19574 96742 19626
rect 96794 19574 96846 19626
rect 96898 19574 118608 19626
rect 1344 19540 118608 19574
rect 1344 18842 118608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 81278 18842
rect 81330 18790 81382 18842
rect 81434 18790 81486 18842
rect 81538 18790 111998 18842
rect 112050 18790 112102 18842
rect 112154 18790 112206 18842
rect 112258 18790 118608 18842
rect 1344 18756 118608 18790
rect 1822 18562 1874 18574
rect 1822 18498 1874 18510
rect 1344 18058 118608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 96638 18058
rect 96690 18006 96742 18058
rect 96794 18006 96846 18058
rect 96898 18006 118608 18058
rect 1344 17972 118608 18006
rect 118078 17554 118130 17566
rect 118078 17490 118130 17502
rect 1822 17442 1874 17454
rect 1822 17378 1874 17390
rect 1344 17274 118608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 81278 17274
rect 81330 17222 81382 17274
rect 81434 17222 81486 17274
rect 81538 17222 111998 17274
rect 112050 17222 112102 17274
rect 112154 17222 112206 17274
rect 112258 17222 118608 17274
rect 1344 17188 118608 17222
rect 118078 16994 118130 17006
rect 118078 16930 118130 16942
rect 1344 16490 118608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 96638 16490
rect 96690 16438 96742 16490
rect 96794 16438 96846 16490
rect 96898 16438 118608 16490
rect 1344 16404 118608 16438
rect 1344 15706 118608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 81278 15706
rect 81330 15654 81382 15706
rect 81434 15654 81486 15706
rect 81538 15654 111998 15706
rect 112050 15654 112102 15706
rect 112154 15654 112206 15706
rect 112258 15654 118608 15706
rect 1344 15620 118608 15654
rect 1344 14922 118608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 96638 14922
rect 96690 14870 96742 14922
rect 96794 14870 96846 14922
rect 96898 14870 118608 14922
rect 1344 14836 118608 14870
rect 118078 14306 118130 14318
rect 118078 14242 118130 14254
rect 1344 14138 118608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 81278 14138
rect 81330 14086 81382 14138
rect 81434 14086 81486 14138
rect 81538 14086 111998 14138
rect 112050 14086 112102 14138
rect 112154 14086 112206 14138
rect 112258 14086 118608 14138
rect 1344 14052 118608 14086
rect 1344 13354 118608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 96638 13354
rect 96690 13302 96742 13354
rect 96794 13302 96846 13354
rect 96898 13302 118608 13354
rect 1344 13268 118608 13302
rect 1344 12570 118608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 81278 12570
rect 81330 12518 81382 12570
rect 81434 12518 81486 12570
rect 81538 12518 111998 12570
rect 112050 12518 112102 12570
rect 112154 12518 112206 12570
rect 112258 12518 118608 12570
rect 1344 12484 118608 12518
rect 118078 12290 118130 12302
rect 118078 12226 118130 12238
rect 1344 11786 118608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 96638 11786
rect 96690 11734 96742 11786
rect 96794 11734 96846 11786
rect 96898 11734 118608 11786
rect 1344 11700 118608 11734
rect 1822 11170 1874 11182
rect 1822 11106 1874 11118
rect 1344 11002 118608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 81278 11002
rect 81330 10950 81382 11002
rect 81434 10950 81486 11002
rect 81538 10950 111998 11002
rect 112050 10950 112102 11002
rect 112154 10950 112206 11002
rect 112258 10950 118608 11002
rect 1344 10916 118608 10950
rect 118078 10722 118130 10734
rect 118078 10658 118130 10670
rect 1344 10218 118608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 96638 10218
rect 96690 10166 96742 10218
rect 96794 10166 96846 10218
rect 96898 10166 118608 10218
rect 1344 10132 118608 10166
rect 1344 9434 118608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 81278 9434
rect 81330 9382 81382 9434
rect 81434 9382 81486 9434
rect 81538 9382 111998 9434
rect 112050 9382 112102 9434
rect 112154 9382 112206 9434
rect 112258 9382 118608 9434
rect 1344 9348 118608 9382
rect 1344 8650 118608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 96638 8650
rect 96690 8598 96742 8650
rect 96794 8598 96846 8650
rect 96898 8598 118608 8650
rect 1344 8564 118608 8598
rect 1822 8034 1874 8046
rect 1822 7970 1874 7982
rect 1344 7866 118608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 81278 7866
rect 81330 7814 81382 7866
rect 81434 7814 81486 7866
rect 81538 7814 111998 7866
rect 112050 7814 112102 7866
rect 112154 7814 112206 7866
rect 112258 7814 118608 7866
rect 1344 7780 118608 7814
rect 1344 7082 118608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 96638 7082
rect 96690 7030 96742 7082
rect 96794 7030 96846 7082
rect 96898 7030 118608 7082
rect 1344 6996 118608 7030
rect 1822 6466 1874 6478
rect 1822 6402 1874 6414
rect 1344 6298 118608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 81278 6298
rect 81330 6246 81382 6298
rect 81434 6246 81486 6298
rect 81538 6246 111998 6298
rect 112050 6246 112102 6298
rect 112154 6246 112206 6298
rect 112258 6246 118608 6298
rect 1344 6212 118608 6246
rect 1344 5514 118608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 96638 5514
rect 96690 5462 96742 5514
rect 96794 5462 96846 5514
rect 96898 5462 118608 5514
rect 1344 5428 118608 5462
rect 1822 4898 1874 4910
rect 1822 4834 1874 4846
rect 118078 4898 118130 4910
rect 118078 4834 118130 4846
rect 1344 4730 118608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 81278 4730
rect 81330 4678 81382 4730
rect 81434 4678 81486 4730
rect 81538 4678 111998 4730
rect 112050 4678 112102 4730
rect 112154 4678 112206 4730
rect 112258 4678 118608 4730
rect 1344 4644 118608 4678
rect 1822 4450 1874 4462
rect 1822 4386 1874 4398
rect 117182 4450 117234 4462
rect 117182 4386 117234 4398
rect 118078 4450 118130 4462
rect 118078 4386 118130 4398
rect 116510 4226 116562 4238
rect 116510 4162 116562 4174
rect 1344 3946 118608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 96638 3946
rect 96690 3894 96742 3946
rect 96794 3894 96846 3946
rect 96898 3894 118608 3946
rect 1344 3860 118608 3894
rect 116834 3502 116846 3554
rect 116898 3502 116910 3554
rect 117730 3390 117742 3442
rect 117794 3390 117806 3442
rect 2270 3330 2322 3342
rect 2270 3266 2322 3278
rect 7646 3330 7698 3342
rect 7646 3266 7698 3278
rect 8318 3330 8370 3342
rect 8318 3266 8370 3278
rect 9662 3330 9714 3342
rect 9662 3266 9714 3278
rect 12350 3330 12402 3342
rect 12350 3266 12402 3278
rect 15038 3330 15090 3342
rect 15038 3266 15090 3278
rect 27134 3330 27186 3342
rect 27134 3266 27186 3278
rect 28366 3330 28418 3342
rect 28366 3266 28418 3278
rect 29822 3330 29874 3342
rect 29822 3266 29874 3278
rect 30494 3330 30546 3342
rect 30494 3266 30546 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 34526 3330 34578 3342
rect 34526 3266 34578 3278
rect 37214 3330 37266 3342
rect 37214 3266 37266 3278
rect 37886 3330 37938 3342
rect 37886 3266 37938 3278
rect 43262 3330 43314 3342
rect 43262 3266 43314 3278
rect 45278 3330 45330 3342
rect 45278 3266 45330 3278
rect 47966 3330 48018 3342
rect 47966 3266 48018 3278
rect 49310 3330 49362 3342
rect 49310 3266 49362 3278
rect 51886 3330 51938 3342
rect 51886 3266 51938 3278
rect 52782 3330 52834 3342
rect 52782 3266 52834 3278
rect 54014 3330 54066 3342
rect 54014 3266 54066 3278
rect 55358 3330 55410 3342
rect 55358 3266 55410 3278
rect 59390 3330 59442 3342
rect 59390 3266 59442 3278
rect 62750 3330 62802 3342
rect 62750 3266 62802 3278
rect 68462 3330 68514 3342
rect 68462 3266 68514 3278
rect 69134 3330 69186 3342
rect 69134 3266 69186 3278
rect 70142 3330 70194 3342
rect 70142 3266 70194 3278
rect 76302 3330 76354 3342
rect 76302 3266 76354 3278
rect 77534 3330 77586 3342
rect 77534 3266 77586 3278
rect 78878 3330 78930 3342
rect 78878 3266 78930 3278
rect 82910 3330 82962 3342
rect 82910 3266 82962 3278
rect 84926 3330 84978 3342
rect 84926 3266 84978 3278
rect 86270 3330 86322 3342
rect 86270 3266 86322 3278
rect 88062 3330 88114 3342
rect 88062 3266 88114 3278
rect 93662 3330 93714 3342
rect 93662 3266 93714 3278
rect 101054 3330 101106 3342
rect 101054 3266 101106 3278
rect 107662 3330 107714 3342
rect 107662 3266 107714 3278
rect 109790 3330 109842 3342
rect 109790 3266 109842 3278
rect 111582 3330 111634 3342
rect 111582 3266 111634 3278
rect 112478 3330 112530 3342
rect 112478 3266 112530 3278
rect 115838 3330 115890 3342
rect 115838 3266 115890 3278
rect 1344 3162 118608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 81278 3162
rect 81330 3110 81382 3162
rect 81434 3110 81486 3162
rect 81538 3110 111998 3162
rect 112050 3110 112102 3162
rect 112154 3110 112206 3162
rect 112258 3110 118608 3162
rect 1344 3076 118608 3110
rect 87378 1822 87390 1874
rect 87442 1871 87454 1874
rect 88050 1871 88062 1874
rect 87442 1825 88062 1871
rect 87442 1822 87454 1825
rect 88050 1822 88062 1825
rect 88114 1822 88126 1874
rect 110898 1822 110910 1874
rect 110962 1871 110974 1874
rect 111570 1871 111582 1874
rect 110962 1825 111582 1871
rect 110962 1822 110974 1825
rect 111570 1822 111582 1825
rect 111634 1822 111646 1874
rect 67890 1710 67902 1762
rect 67954 1759 67966 1762
rect 68450 1759 68462 1762
rect 67954 1713 68462 1759
rect 67954 1710 67966 1713
rect 68450 1710 68462 1713
rect 68514 1710 68526 1762
<< via1 >>
rect 60510 132638 60562 132690
rect 61518 132638 61570 132690
rect 102846 132638 102898 132690
rect 103742 132638 103794 132690
rect 4478 132470 4530 132522
rect 4582 132470 4634 132522
rect 4686 132470 4738 132522
rect 35198 132470 35250 132522
rect 35302 132470 35354 132522
rect 35406 132470 35458 132522
rect 65918 132470 65970 132522
rect 66022 132470 66074 132522
rect 66126 132470 66178 132522
rect 96638 132470 96690 132522
rect 96742 132470 96794 132522
rect 96846 132470 96898 132522
rect 22094 132190 22146 132242
rect 59838 132190 59890 132242
rect 21422 132078 21474 132130
rect 60846 132078 60898 132130
rect 1822 131966 1874 132018
rect 2494 131966 2546 132018
rect 10334 131966 10386 132018
rect 11678 131966 11730 132018
rect 13582 131966 13634 132018
rect 23774 131966 23826 132018
rect 26462 131966 26514 132018
rect 27806 131966 27858 132018
rect 29822 131966 29874 132018
rect 31166 131966 31218 132018
rect 36318 131966 36370 132018
rect 37214 131966 37266 132018
rect 39902 131966 39954 132018
rect 45950 131966 46002 132018
rect 51326 131966 51378 132018
rect 53342 131966 53394 132018
rect 54686 131966 54738 132018
rect 58718 131966 58770 132018
rect 61518 131966 61570 132018
rect 63422 131966 63474 132018
rect 64766 131966 64818 132018
rect 66110 131966 66162 132018
rect 67454 131966 67506 132018
rect 69470 131966 69522 132018
rect 72382 131966 72434 132018
rect 73502 131966 73554 132018
rect 74846 131966 74898 132018
rect 76302 131966 76354 132018
rect 80894 131966 80946 132018
rect 82238 131966 82290 132018
rect 84254 131966 84306 132018
rect 85598 131966 85650 132018
rect 88286 131966 88338 132018
rect 89630 131966 89682 132018
rect 95902 131966 95954 132018
rect 103742 131966 103794 132018
rect 104414 131966 104466 132018
rect 109118 131966 109170 132018
rect 115502 131966 115554 132018
rect 116510 131966 116562 132018
rect 117294 131966 117346 132018
rect 117854 131966 117906 132018
rect 20638 131854 20690 131906
rect 60622 131854 60674 131906
rect 19838 131686 19890 131738
rect 19942 131686 19994 131738
rect 20046 131686 20098 131738
rect 50558 131686 50610 131738
rect 50662 131686 50714 131738
rect 50766 131686 50818 131738
rect 81278 131686 81330 131738
rect 81382 131686 81434 131738
rect 81486 131686 81538 131738
rect 111998 131686 112050 131738
rect 112102 131686 112154 131738
rect 112206 131686 112258 131738
rect 4478 130902 4530 130954
rect 4582 130902 4634 130954
rect 4686 130902 4738 130954
rect 35198 130902 35250 130954
rect 35302 130902 35354 130954
rect 35406 130902 35458 130954
rect 65918 130902 65970 130954
rect 66022 130902 66074 130954
rect 66126 130902 66178 130954
rect 96638 130902 96690 130954
rect 96742 130902 96794 130954
rect 96846 130902 96898 130954
rect 1822 130398 1874 130450
rect 19838 130118 19890 130170
rect 19942 130118 19994 130170
rect 20046 130118 20098 130170
rect 50558 130118 50610 130170
rect 50662 130118 50714 130170
rect 50766 130118 50818 130170
rect 81278 130118 81330 130170
rect 81382 130118 81434 130170
rect 81486 130118 81538 130170
rect 111998 130118 112050 130170
rect 112102 130118 112154 130170
rect 112206 130118 112258 130170
rect 4478 129334 4530 129386
rect 4582 129334 4634 129386
rect 4686 129334 4738 129386
rect 35198 129334 35250 129386
rect 35302 129334 35354 129386
rect 35406 129334 35458 129386
rect 65918 129334 65970 129386
rect 66022 129334 66074 129386
rect 66126 129334 66178 129386
rect 96638 129334 96690 129386
rect 96742 129334 96794 129386
rect 96846 129334 96898 129386
rect 19838 128550 19890 128602
rect 19942 128550 19994 128602
rect 20046 128550 20098 128602
rect 50558 128550 50610 128602
rect 50662 128550 50714 128602
rect 50766 128550 50818 128602
rect 81278 128550 81330 128602
rect 81382 128550 81434 128602
rect 81486 128550 81538 128602
rect 111998 128550 112050 128602
rect 112102 128550 112154 128602
rect 112206 128550 112258 128602
rect 1822 128270 1874 128322
rect 4478 127766 4530 127818
rect 4582 127766 4634 127818
rect 4686 127766 4738 127818
rect 35198 127766 35250 127818
rect 35302 127766 35354 127818
rect 35406 127766 35458 127818
rect 65918 127766 65970 127818
rect 66022 127766 66074 127818
rect 66126 127766 66178 127818
rect 96638 127766 96690 127818
rect 96742 127766 96794 127818
rect 96846 127766 96898 127818
rect 1822 127150 1874 127202
rect 19838 126982 19890 127034
rect 19942 126982 19994 127034
rect 20046 126982 20098 127034
rect 50558 126982 50610 127034
rect 50662 126982 50714 127034
rect 50766 126982 50818 127034
rect 81278 126982 81330 127034
rect 81382 126982 81434 127034
rect 81486 126982 81538 127034
rect 111998 126982 112050 127034
rect 112102 126982 112154 127034
rect 112206 126982 112258 127034
rect 118078 126702 118130 126754
rect 4478 126198 4530 126250
rect 4582 126198 4634 126250
rect 4686 126198 4738 126250
rect 35198 126198 35250 126250
rect 35302 126198 35354 126250
rect 35406 126198 35458 126250
rect 65918 126198 65970 126250
rect 66022 126198 66074 126250
rect 66126 126198 66178 126250
rect 96638 126198 96690 126250
rect 96742 126198 96794 126250
rect 96846 126198 96898 126250
rect 19838 125414 19890 125466
rect 19942 125414 19994 125466
rect 20046 125414 20098 125466
rect 50558 125414 50610 125466
rect 50662 125414 50714 125466
rect 50766 125414 50818 125466
rect 81278 125414 81330 125466
rect 81382 125414 81434 125466
rect 81486 125414 81538 125466
rect 111998 125414 112050 125466
rect 112102 125414 112154 125466
rect 112206 125414 112258 125466
rect 1822 125134 1874 125186
rect 4478 124630 4530 124682
rect 4582 124630 4634 124682
rect 4686 124630 4738 124682
rect 35198 124630 35250 124682
rect 35302 124630 35354 124682
rect 35406 124630 35458 124682
rect 65918 124630 65970 124682
rect 66022 124630 66074 124682
rect 66126 124630 66178 124682
rect 96638 124630 96690 124682
rect 96742 124630 96794 124682
rect 96846 124630 96898 124682
rect 118078 124014 118130 124066
rect 19838 123846 19890 123898
rect 19942 123846 19994 123898
rect 20046 123846 20098 123898
rect 50558 123846 50610 123898
rect 50662 123846 50714 123898
rect 50766 123846 50818 123898
rect 81278 123846 81330 123898
rect 81382 123846 81434 123898
rect 81486 123846 81538 123898
rect 111998 123846 112050 123898
rect 112102 123846 112154 123898
rect 112206 123846 112258 123898
rect 1822 123566 1874 123618
rect 4478 123062 4530 123114
rect 4582 123062 4634 123114
rect 4686 123062 4738 123114
rect 35198 123062 35250 123114
rect 35302 123062 35354 123114
rect 35406 123062 35458 123114
rect 65918 123062 65970 123114
rect 66022 123062 66074 123114
rect 66126 123062 66178 123114
rect 96638 123062 96690 123114
rect 96742 123062 96794 123114
rect 96846 123062 96898 123114
rect 19838 122278 19890 122330
rect 19942 122278 19994 122330
rect 20046 122278 20098 122330
rect 50558 122278 50610 122330
rect 50662 122278 50714 122330
rect 50766 122278 50818 122330
rect 81278 122278 81330 122330
rect 81382 122278 81434 122330
rect 81486 122278 81538 122330
rect 111998 122278 112050 122330
rect 112102 122278 112154 122330
rect 112206 122278 112258 122330
rect 1822 121998 1874 122050
rect 4478 121494 4530 121546
rect 4582 121494 4634 121546
rect 4686 121494 4738 121546
rect 35198 121494 35250 121546
rect 35302 121494 35354 121546
rect 35406 121494 35458 121546
rect 65918 121494 65970 121546
rect 66022 121494 66074 121546
rect 66126 121494 66178 121546
rect 96638 121494 96690 121546
rect 96742 121494 96794 121546
rect 96846 121494 96898 121546
rect 19838 120710 19890 120762
rect 19942 120710 19994 120762
rect 20046 120710 20098 120762
rect 50558 120710 50610 120762
rect 50662 120710 50714 120762
rect 50766 120710 50818 120762
rect 81278 120710 81330 120762
rect 81382 120710 81434 120762
rect 81486 120710 81538 120762
rect 111998 120710 112050 120762
rect 112102 120710 112154 120762
rect 112206 120710 112258 120762
rect 4478 119926 4530 119978
rect 4582 119926 4634 119978
rect 4686 119926 4738 119978
rect 35198 119926 35250 119978
rect 35302 119926 35354 119978
rect 35406 119926 35458 119978
rect 65918 119926 65970 119978
rect 66022 119926 66074 119978
rect 66126 119926 66178 119978
rect 96638 119926 96690 119978
rect 96742 119926 96794 119978
rect 96846 119926 96898 119978
rect 19838 119142 19890 119194
rect 19942 119142 19994 119194
rect 20046 119142 20098 119194
rect 50558 119142 50610 119194
rect 50662 119142 50714 119194
rect 50766 119142 50818 119194
rect 81278 119142 81330 119194
rect 81382 119142 81434 119194
rect 81486 119142 81538 119194
rect 111998 119142 112050 119194
rect 112102 119142 112154 119194
rect 112206 119142 112258 119194
rect 4478 118358 4530 118410
rect 4582 118358 4634 118410
rect 4686 118358 4738 118410
rect 35198 118358 35250 118410
rect 35302 118358 35354 118410
rect 35406 118358 35458 118410
rect 65918 118358 65970 118410
rect 66022 118358 66074 118410
rect 66126 118358 66178 118410
rect 96638 118358 96690 118410
rect 96742 118358 96794 118410
rect 96846 118358 96898 118410
rect 19838 117574 19890 117626
rect 19942 117574 19994 117626
rect 20046 117574 20098 117626
rect 50558 117574 50610 117626
rect 50662 117574 50714 117626
rect 50766 117574 50818 117626
rect 81278 117574 81330 117626
rect 81382 117574 81434 117626
rect 81486 117574 81538 117626
rect 111998 117574 112050 117626
rect 112102 117574 112154 117626
rect 112206 117574 112258 117626
rect 1822 117294 1874 117346
rect 4478 116790 4530 116842
rect 4582 116790 4634 116842
rect 4686 116790 4738 116842
rect 35198 116790 35250 116842
rect 35302 116790 35354 116842
rect 35406 116790 35458 116842
rect 65918 116790 65970 116842
rect 66022 116790 66074 116842
rect 66126 116790 66178 116842
rect 96638 116790 96690 116842
rect 96742 116790 96794 116842
rect 96846 116790 96898 116842
rect 118078 116286 118130 116338
rect 19838 116006 19890 116058
rect 19942 116006 19994 116058
rect 20046 116006 20098 116058
rect 50558 116006 50610 116058
rect 50662 116006 50714 116058
rect 50766 116006 50818 116058
rect 81278 116006 81330 116058
rect 81382 116006 81434 116058
rect 81486 116006 81538 116058
rect 111998 116006 112050 116058
rect 112102 116006 112154 116058
rect 112206 116006 112258 116058
rect 118078 115726 118130 115778
rect 4478 115222 4530 115274
rect 4582 115222 4634 115274
rect 4686 115222 4738 115274
rect 35198 115222 35250 115274
rect 35302 115222 35354 115274
rect 35406 115222 35458 115274
rect 65918 115222 65970 115274
rect 66022 115222 66074 115274
rect 66126 115222 66178 115274
rect 96638 115222 96690 115274
rect 96742 115222 96794 115274
rect 96846 115222 96898 115274
rect 19838 114438 19890 114490
rect 19942 114438 19994 114490
rect 20046 114438 20098 114490
rect 50558 114438 50610 114490
rect 50662 114438 50714 114490
rect 50766 114438 50818 114490
rect 81278 114438 81330 114490
rect 81382 114438 81434 114490
rect 81486 114438 81538 114490
rect 111998 114438 112050 114490
rect 112102 114438 112154 114490
rect 112206 114438 112258 114490
rect 118078 114270 118130 114322
rect 4478 113654 4530 113706
rect 4582 113654 4634 113706
rect 4686 113654 4738 113706
rect 35198 113654 35250 113706
rect 35302 113654 35354 113706
rect 35406 113654 35458 113706
rect 65918 113654 65970 113706
rect 66022 113654 66074 113706
rect 66126 113654 66178 113706
rect 96638 113654 96690 113706
rect 96742 113654 96794 113706
rect 96846 113654 96898 113706
rect 19838 112870 19890 112922
rect 19942 112870 19994 112922
rect 20046 112870 20098 112922
rect 50558 112870 50610 112922
rect 50662 112870 50714 112922
rect 50766 112870 50818 112922
rect 81278 112870 81330 112922
rect 81382 112870 81434 112922
rect 81486 112870 81538 112922
rect 111998 112870 112050 112922
rect 112102 112870 112154 112922
rect 112206 112870 112258 112922
rect 4478 112086 4530 112138
rect 4582 112086 4634 112138
rect 4686 112086 4738 112138
rect 35198 112086 35250 112138
rect 35302 112086 35354 112138
rect 35406 112086 35458 112138
rect 65918 112086 65970 112138
rect 66022 112086 66074 112138
rect 66126 112086 66178 112138
rect 96638 112086 96690 112138
rect 96742 112086 96794 112138
rect 96846 112086 96898 112138
rect 118078 111582 118130 111634
rect 1822 111470 1874 111522
rect 19838 111302 19890 111354
rect 19942 111302 19994 111354
rect 20046 111302 20098 111354
rect 50558 111302 50610 111354
rect 50662 111302 50714 111354
rect 50766 111302 50818 111354
rect 81278 111302 81330 111354
rect 81382 111302 81434 111354
rect 81486 111302 81538 111354
rect 111998 111302 112050 111354
rect 112102 111302 112154 111354
rect 112206 111302 112258 111354
rect 118078 111022 118130 111074
rect 4478 110518 4530 110570
rect 4582 110518 4634 110570
rect 4686 110518 4738 110570
rect 35198 110518 35250 110570
rect 35302 110518 35354 110570
rect 35406 110518 35458 110570
rect 65918 110518 65970 110570
rect 66022 110518 66074 110570
rect 66126 110518 66178 110570
rect 96638 110518 96690 110570
rect 96742 110518 96794 110570
rect 96846 110518 96898 110570
rect 1822 109902 1874 109954
rect 19838 109734 19890 109786
rect 19942 109734 19994 109786
rect 20046 109734 20098 109786
rect 50558 109734 50610 109786
rect 50662 109734 50714 109786
rect 50766 109734 50818 109786
rect 81278 109734 81330 109786
rect 81382 109734 81434 109786
rect 81486 109734 81538 109786
rect 111998 109734 112050 109786
rect 112102 109734 112154 109786
rect 112206 109734 112258 109786
rect 4478 108950 4530 109002
rect 4582 108950 4634 109002
rect 4686 108950 4738 109002
rect 35198 108950 35250 109002
rect 35302 108950 35354 109002
rect 35406 108950 35458 109002
rect 65918 108950 65970 109002
rect 66022 108950 66074 109002
rect 66126 108950 66178 109002
rect 96638 108950 96690 109002
rect 96742 108950 96794 109002
rect 96846 108950 96898 109002
rect 19838 108166 19890 108218
rect 19942 108166 19994 108218
rect 20046 108166 20098 108218
rect 50558 108166 50610 108218
rect 50662 108166 50714 108218
rect 50766 108166 50818 108218
rect 81278 108166 81330 108218
rect 81382 108166 81434 108218
rect 81486 108166 81538 108218
rect 111998 108166 112050 108218
rect 112102 108166 112154 108218
rect 112206 108166 112258 108218
rect 118078 107886 118130 107938
rect 4478 107382 4530 107434
rect 4582 107382 4634 107434
rect 4686 107382 4738 107434
rect 35198 107382 35250 107434
rect 35302 107382 35354 107434
rect 35406 107382 35458 107434
rect 65918 107382 65970 107434
rect 66022 107382 66074 107434
rect 66126 107382 66178 107434
rect 96638 107382 96690 107434
rect 96742 107382 96794 107434
rect 96846 107382 96898 107434
rect 118078 106766 118130 106818
rect 19838 106598 19890 106650
rect 19942 106598 19994 106650
rect 20046 106598 20098 106650
rect 50558 106598 50610 106650
rect 50662 106598 50714 106650
rect 50766 106598 50818 106650
rect 81278 106598 81330 106650
rect 81382 106598 81434 106650
rect 81486 106598 81538 106650
rect 111998 106598 112050 106650
rect 112102 106598 112154 106650
rect 112206 106598 112258 106650
rect 4478 105814 4530 105866
rect 4582 105814 4634 105866
rect 4686 105814 4738 105866
rect 35198 105814 35250 105866
rect 35302 105814 35354 105866
rect 35406 105814 35458 105866
rect 65918 105814 65970 105866
rect 66022 105814 66074 105866
rect 66126 105814 66178 105866
rect 96638 105814 96690 105866
rect 96742 105814 96794 105866
rect 96846 105814 96898 105866
rect 1822 105198 1874 105250
rect 19838 105030 19890 105082
rect 19942 105030 19994 105082
rect 20046 105030 20098 105082
rect 50558 105030 50610 105082
rect 50662 105030 50714 105082
rect 50766 105030 50818 105082
rect 81278 105030 81330 105082
rect 81382 105030 81434 105082
rect 81486 105030 81538 105082
rect 111998 105030 112050 105082
rect 112102 105030 112154 105082
rect 112206 105030 112258 105082
rect 4478 104246 4530 104298
rect 4582 104246 4634 104298
rect 4686 104246 4738 104298
rect 35198 104246 35250 104298
rect 35302 104246 35354 104298
rect 35406 104246 35458 104298
rect 65918 104246 65970 104298
rect 66022 104246 66074 104298
rect 66126 104246 66178 104298
rect 96638 104246 96690 104298
rect 96742 104246 96794 104298
rect 96846 104246 96898 104298
rect 19838 103462 19890 103514
rect 19942 103462 19994 103514
rect 20046 103462 20098 103514
rect 50558 103462 50610 103514
rect 50662 103462 50714 103514
rect 50766 103462 50818 103514
rect 81278 103462 81330 103514
rect 81382 103462 81434 103514
rect 81486 103462 81538 103514
rect 111998 103462 112050 103514
rect 112102 103462 112154 103514
rect 112206 103462 112258 103514
rect 118078 103182 118130 103234
rect 4478 102678 4530 102730
rect 4582 102678 4634 102730
rect 4686 102678 4738 102730
rect 35198 102678 35250 102730
rect 35302 102678 35354 102730
rect 35406 102678 35458 102730
rect 65918 102678 65970 102730
rect 66022 102678 66074 102730
rect 66126 102678 66178 102730
rect 96638 102678 96690 102730
rect 96742 102678 96794 102730
rect 96846 102678 96898 102730
rect 19838 101894 19890 101946
rect 19942 101894 19994 101946
rect 20046 101894 20098 101946
rect 50558 101894 50610 101946
rect 50662 101894 50714 101946
rect 50766 101894 50818 101946
rect 81278 101894 81330 101946
rect 81382 101894 81434 101946
rect 81486 101894 81538 101946
rect 111998 101894 112050 101946
rect 112102 101894 112154 101946
rect 112206 101894 112258 101946
rect 1822 101614 1874 101666
rect 4478 101110 4530 101162
rect 4582 101110 4634 101162
rect 4686 101110 4738 101162
rect 35198 101110 35250 101162
rect 35302 101110 35354 101162
rect 35406 101110 35458 101162
rect 65918 101110 65970 101162
rect 66022 101110 66074 101162
rect 66126 101110 66178 101162
rect 96638 101110 96690 101162
rect 96742 101110 96794 101162
rect 96846 101110 96898 101162
rect 19838 100326 19890 100378
rect 19942 100326 19994 100378
rect 20046 100326 20098 100378
rect 50558 100326 50610 100378
rect 50662 100326 50714 100378
rect 50766 100326 50818 100378
rect 81278 100326 81330 100378
rect 81382 100326 81434 100378
rect 81486 100326 81538 100378
rect 111998 100326 112050 100378
rect 112102 100326 112154 100378
rect 112206 100326 112258 100378
rect 4478 99542 4530 99594
rect 4582 99542 4634 99594
rect 4686 99542 4738 99594
rect 35198 99542 35250 99594
rect 35302 99542 35354 99594
rect 35406 99542 35458 99594
rect 65918 99542 65970 99594
rect 66022 99542 66074 99594
rect 66126 99542 66178 99594
rect 96638 99542 96690 99594
rect 96742 99542 96794 99594
rect 96846 99542 96898 99594
rect 19838 98758 19890 98810
rect 19942 98758 19994 98810
rect 20046 98758 20098 98810
rect 50558 98758 50610 98810
rect 50662 98758 50714 98810
rect 50766 98758 50818 98810
rect 81278 98758 81330 98810
rect 81382 98758 81434 98810
rect 81486 98758 81538 98810
rect 111998 98758 112050 98810
rect 112102 98758 112154 98810
rect 112206 98758 112258 98810
rect 118078 98478 118130 98530
rect 4478 97974 4530 98026
rect 4582 97974 4634 98026
rect 4686 97974 4738 98026
rect 35198 97974 35250 98026
rect 35302 97974 35354 98026
rect 35406 97974 35458 98026
rect 65918 97974 65970 98026
rect 66022 97974 66074 98026
rect 66126 97974 66178 98026
rect 96638 97974 96690 98026
rect 96742 97974 96794 98026
rect 96846 97974 96898 98026
rect 118078 97358 118130 97410
rect 19838 97190 19890 97242
rect 19942 97190 19994 97242
rect 20046 97190 20098 97242
rect 50558 97190 50610 97242
rect 50662 97190 50714 97242
rect 50766 97190 50818 97242
rect 81278 97190 81330 97242
rect 81382 97190 81434 97242
rect 81486 97190 81538 97242
rect 111998 97190 112050 97242
rect 112102 97190 112154 97242
rect 112206 97190 112258 97242
rect 1822 96910 1874 96962
rect 4478 96406 4530 96458
rect 4582 96406 4634 96458
rect 4686 96406 4738 96458
rect 35198 96406 35250 96458
rect 35302 96406 35354 96458
rect 35406 96406 35458 96458
rect 65918 96406 65970 96458
rect 66022 96406 66074 96458
rect 66126 96406 66178 96458
rect 96638 96406 96690 96458
rect 96742 96406 96794 96458
rect 96846 96406 96898 96458
rect 118078 95790 118130 95842
rect 19838 95622 19890 95674
rect 19942 95622 19994 95674
rect 20046 95622 20098 95674
rect 50558 95622 50610 95674
rect 50662 95622 50714 95674
rect 50766 95622 50818 95674
rect 81278 95622 81330 95674
rect 81382 95622 81434 95674
rect 81486 95622 81538 95674
rect 111998 95622 112050 95674
rect 112102 95622 112154 95674
rect 112206 95622 112258 95674
rect 1822 95342 1874 95394
rect 4478 94838 4530 94890
rect 4582 94838 4634 94890
rect 4686 94838 4738 94890
rect 35198 94838 35250 94890
rect 35302 94838 35354 94890
rect 35406 94838 35458 94890
rect 65918 94838 65970 94890
rect 66022 94838 66074 94890
rect 66126 94838 66178 94890
rect 96638 94838 96690 94890
rect 96742 94838 96794 94890
rect 96846 94838 96898 94890
rect 19838 94054 19890 94106
rect 19942 94054 19994 94106
rect 20046 94054 20098 94106
rect 50558 94054 50610 94106
rect 50662 94054 50714 94106
rect 50766 94054 50818 94106
rect 81278 94054 81330 94106
rect 81382 94054 81434 94106
rect 81486 94054 81538 94106
rect 111998 94054 112050 94106
rect 112102 94054 112154 94106
rect 112206 94054 112258 94106
rect 4478 93270 4530 93322
rect 4582 93270 4634 93322
rect 4686 93270 4738 93322
rect 35198 93270 35250 93322
rect 35302 93270 35354 93322
rect 35406 93270 35458 93322
rect 65918 93270 65970 93322
rect 66022 93270 66074 93322
rect 66126 93270 66178 93322
rect 96638 93270 96690 93322
rect 96742 93270 96794 93322
rect 96846 93270 96898 93322
rect 1822 92654 1874 92706
rect 19838 92486 19890 92538
rect 19942 92486 19994 92538
rect 20046 92486 20098 92538
rect 50558 92486 50610 92538
rect 50662 92486 50714 92538
rect 50766 92486 50818 92538
rect 81278 92486 81330 92538
rect 81382 92486 81434 92538
rect 81486 92486 81538 92538
rect 111998 92486 112050 92538
rect 112102 92486 112154 92538
rect 112206 92486 112258 92538
rect 4478 91702 4530 91754
rect 4582 91702 4634 91754
rect 4686 91702 4738 91754
rect 35198 91702 35250 91754
rect 35302 91702 35354 91754
rect 35406 91702 35458 91754
rect 65918 91702 65970 91754
rect 66022 91702 66074 91754
rect 66126 91702 66178 91754
rect 96638 91702 96690 91754
rect 96742 91702 96794 91754
rect 96846 91702 96898 91754
rect 1822 91086 1874 91138
rect 118078 91086 118130 91138
rect 19838 90918 19890 90970
rect 19942 90918 19994 90970
rect 20046 90918 20098 90970
rect 50558 90918 50610 90970
rect 50662 90918 50714 90970
rect 50766 90918 50818 90970
rect 81278 90918 81330 90970
rect 81382 90918 81434 90970
rect 81486 90918 81538 90970
rect 111998 90918 112050 90970
rect 112102 90918 112154 90970
rect 112206 90918 112258 90970
rect 2158 90638 2210 90690
rect 1822 90526 1874 90578
rect 4478 90134 4530 90186
rect 4582 90134 4634 90186
rect 4686 90134 4738 90186
rect 35198 90134 35250 90186
rect 35302 90134 35354 90186
rect 35406 90134 35458 90186
rect 65918 90134 65970 90186
rect 66022 90134 66074 90186
rect 66126 90134 66178 90186
rect 96638 90134 96690 90186
rect 96742 90134 96794 90186
rect 96846 90134 96898 90186
rect 1822 89854 1874 89906
rect 19838 89350 19890 89402
rect 19942 89350 19994 89402
rect 20046 89350 20098 89402
rect 50558 89350 50610 89402
rect 50662 89350 50714 89402
rect 50766 89350 50818 89402
rect 81278 89350 81330 89402
rect 81382 89350 81434 89402
rect 81486 89350 81538 89402
rect 111998 89350 112050 89402
rect 112102 89350 112154 89402
rect 112206 89350 112258 89402
rect 4478 88566 4530 88618
rect 4582 88566 4634 88618
rect 4686 88566 4738 88618
rect 35198 88566 35250 88618
rect 35302 88566 35354 88618
rect 35406 88566 35458 88618
rect 65918 88566 65970 88618
rect 66022 88566 66074 88618
rect 66126 88566 66178 88618
rect 96638 88566 96690 88618
rect 96742 88566 96794 88618
rect 96846 88566 96898 88618
rect 118078 88062 118130 88114
rect 19838 87782 19890 87834
rect 19942 87782 19994 87834
rect 20046 87782 20098 87834
rect 50558 87782 50610 87834
rect 50662 87782 50714 87834
rect 50766 87782 50818 87834
rect 81278 87782 81330 87834
rect 81382 87782 81434 87834
rect 81486 87782 81538 87834
rect 111998 87782 112050 87834
rect 112102 87782 112154 87834
rect 112206 87782 112258 87834
rect 4478 86998 4530 87050
rect 4582 86998 4634 87050
rect 4686 86998 4738 87050
rect 35198 86998 35250 87050
rect 35302 86998 35354 87050
rect 35406 86998 35458 87050
rect 65918 86998 65970 87050
rect 66022 86998 66074 87050
rect 66126 86998 66178 87050
rect 96638 86998 96690 87050
rect 96742 86998 96794 87050
rect 96846 86998 96898 87050
rect 19838 86214 19890 86266
rect 19942 86214 19994 86266
rect 20046 86214 20098 86266
rect 50558 86214 50610 86266
rect 50662 86214 50714 86266
rect 50766 86214 50818 86266
rect 81278 86214 81330 86266
rect 81382 86214 81434 86266
rect 81486 86214 81538 86266
rect 111998 86214 112050 86266
rect 112102 86214 112154 86266
rect 112206 86214 112258 86266
rect 4478 85430 4530 85482
rect 4582 85430 4634 85482
rect 4686 85430 4738 85482
rect 35198 85430 35250 85482
rect 35302 85430 35354 85482
rect 35406 85430 35458 85482
rect 65918 85430 65970 85482
rect 66022 85430 66074 85482
rect 66126 85430 66178 85482
rect 96638 85430 96690 85482
rect 96742 85430 96794 85482
rect 96846 85430 96898 85482
rect 2830 85038 2882 85090
rect 2158 84926 2210 84978
rect 3502 84814 3554 84866
rect 19838 84646 19890 84698
rect 19942 84646 19994 84698
rect 20046 84646 20098 84698
rect 50558 84646 50610 84698
rect 50662 84646 50714 84698
rect 50766 84646 50818 84698
rect 81278 84646 81330 84698
rect 81382 84646 81434 84698
rect 81486 84646 81538 84698
rect 111998 84646 112050 84698
rect 112102 84646 112154 84698
rect 112206 84646 112258 84698
rect 118078 84366 118130 84418
rect 4478 83862 4530 83914
rect 4582 83862 4634 83914
rect 4686 83862 4738 83914
rect 35198 83862 35250 83914
rect 35302 83862 35354 83914
rect 35406 83862 35458 83914
rect 65918 83862 65970 83914
rect 66022 83862 66074 83914
rect 66126 83862 66178 83914
rect 96638 83862 96690 83914
rect 96742 83862 96794 83914
rect 96846 83862 96898 83914
rect 2494 83358 2546 83410
rect 1822 83246 1874 83298
rect 19838 83078 19890 83130
rect 19942 83078 19994 83130
rect 20046 83078 20098 83130
rect 50558 83078 50610 83130
rect 50662 83078 50714 83130
rect 50766 83078 50818 83130
rect 81278 83078 81330 83130
rect 81382 83078 81434 83130
rect 81486 83078 81538 83130
rect 111998 83078 112050 83130
rect 112102 83078 112154 83130
rect 112206 83078 112258 83130
rect 118078 82798 118130 82850
rect 4478 82294 4530 82346
rect 4582 82294 4634 82346
rect 4686 82294 4738 82346
rect 35198 82294 35250 82346
rect 35302 82294 35354 82346
rect 35406 82294 35458 82346
rect 65918 82294 65970 82346
rect 66022 82294 66074 82346
rect 66126 82294 66178 82346
rect 96638 82294 96690 82346
rect 96742 82294 96794 82346
rect 96846 82294 96898 82346
rect 19838 81510 19890 81562
rect 19942 81510 19994 81562
rect 20046 81510 20098 81562
rect 50558 81510 50610 81562
rect 50662 81510 50714 81562
rect 50766 81510 50818 81562
rect 81278 81510 81330 81562
rect 81382 81510 81434 81562
rect 81486 81510 81538 81562
rect 111998 81510 112050 81562
rect 112102 81510 112154 81562
rect 112206 81510 112258 81562
rect 4478 80726 4530 80778
rect 4582 80726 4634 80778
rect 4686 80726 4738 80778
rect 35198 80726 35250 80778
rect 35302 80726 35354 80778
rect 35406 80726 35458 80778
rect 65918 80726 65970 80778
rect 66022 80726 66074 80778
rect 66126 80726 66178 80778
rect 96638 80726 96690 80778
rect 96742 80726 96794 80778
rect 96846 80726 96898 80778
rect 19838 79942 19890 79994
rect 19942 79942 19994 79994
rect 20046 79942 20098 79994
rect 50558 79942 50610 79994
rect 50662 79942 50714 79994
rect 50766 79942 50818 79994
rect 81278 79942 81330 79994
rect 81382 79942 81434 79994
rect 81486 79942 81538 79994
rect 111998 79942 112050 79994
rect 112102 79942 112154 79994
rect 112206 79942 112258 79994
rect 118078 79662 118130 79714
rect 4478 79158 4530 79210
rect 4582 79158 4634 79210
rect 4686 79158 4738 79210
rect 35198 79158 35250 79210
rect 35302 79158 35354 79210
rect 35406 79158 35458 79210
rect 65918 79158 65970 79210
rect 66022 79158 66074 79210
rect 66126 79158 66178 79210
rect 96638 79158 96690 79210
rect 96742 79158 96794 79210
rect 96846 79158 96898 79210
rect 19838 78374 19890 78426
rect 19942 78374 19994 78426
rect 20046 78374 20098 78426
rect 50558 78374 50610 78426
rect 50662 78374 50714 78426
rect 50766 78374 50818 78426
rect 81278 78374 81330 78426
rect 81382 78374 81434 78426
rect 81486 78374 81538 78426
rect 111998 78374 112050 78426
rect 112102 78374 112154 78426
rect 112206 78374 112258 78426
rect 2158 78094 2210 78146
rect 1822 77982 1874 78034
rect 4478 77590 4530 77642
rect 4582 77590 4634 77642
rect 4686 77590 4738 77642
rect 35198 77590 35250 77642
rect 35302 77590 35354 77642
rect 35406 77590 35458 77642
rect 65918 77590 65970 77642
rect 66022 77590 66074 77642
rect 66126 77590 66178 77642
rect 96638 77590 96690 77642
rect 96742 77590 96794 77642
rect 96846 77590 96898 77642
rect 1822 77310 1874 77362
rect 118078 76974 118130 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 81278 76806 81330 76858
rect 81382 76806 81434 76858
rect 81486 76806 81538 76858
rect 111998 76806 112050 76858
rect 112102 76806 112154 76858
rect 112206 76806 112258 76858
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 96638 76022 96690 76074
rect 96742 76022 96794 76074
rect 96846 76022 96898 76074
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 81278 75238 81330 75290
rect 81382 75238 81434 75290
rect 81486 75238 81538 75290
rect 111998 75238 112050 75290
rect 112102 75238 112154 75290
rect 112206 75238 112258 75290
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 96638 74454 96690 74506
rect 96742 74454 96794 74506
rect 96846 74454 96898 74506
rect 118078 73838 118130 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 81278 73670 81330 73722
rect 81382 73670 81434 73722
rect 81486 73670 81538 73722
rect 111998 73670 112050 73722
rect 112102 73670 112154 73722
rect 112206 73670 112258 73722
rect 1822 73390 1874 73442
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 96638 72886 96690 72938
rect 96742 72886 96794 72938
rect 96846 72886 96898 72938
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 81278 72102 81330 72154
rect 81382 72102 81434 72154
rect 81486 72102 81538 72154
rect 111998 72102 112050 72154
rect 112102 72102 112154 72154
rect 112206 72102 112258 72154
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 96638 71318 96690 71370
rect 96742 71318 96794 71370
rect 96846 71318 96898 71370
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 81278 70534 81330 70586
rect 81382 70534 81434 70586
rect 81486 70534 81538 70586
rect 111998 70534 112050 70586
rect 112102 70534 112154 70586
rect 112206 70534 112258 70586
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 96638 69750 96690 69802
rect 96742 69750 96794 69802
rect 96846 69750 96898 69802
rect 118078 69246 118130 69298
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 81278 68966 81330 69018
rect 81382 68966 81434 69018
rect 81486 68966 81538 69018
rect 111998 68966 112050 69018
rect 112102 68966 112154 69018
rect 112206 68966 112258 69018
rect 3166 68798 3218 68850
rect 20078 68798 20130 68850
rect 2606 68686 2658 68738
rect 118078 68686 118130 68738
rect 19966 68462 20018 68514
rect 20638 68462 20690 68514
rect 2718 68350 2770 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 96638 68182 96690 68234
rect 96742 68182 96794 68234
rect 96846 68182 96898 68234
rect 60062 67902 60114 67954
rect 3390 67790 3442 67842
rect 4062 67790 4114 67842
rect 59614 67790 59666 67842
rect 2046 67678 2098 67730
rect 2494 67678 2546 67730
rect 2830 67678 2882 67730
rect 3502 67566 3554 67618
rect 3726 67566 3778 67618
rect 59278 67566 59330 67618
rect 118078 67566 118130 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 81278 67398 81330 67450
rect 81382 67398 81434 67450
rect 81486 67398 81538 67450
rect 111998 67398 112050 67450
rect 112102 67398 112154 67450
rect 112206 67398 112258 67450
rect 6302 67118 6354 67170
rect 1934 67006 1986 67058
rect 2270 67006 2322 67058
rect 4622 67006 4674 67058
rect 5070 67006 5122 67058
rect 5854 66782 5906 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 96638 66614 96690 66666
rect 96742 66614 96794 66666
rect 96846 66614 96898 66666
rect 1822 66222 1874 66274
rect 2158 66110 2210 66162
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 81278 65830 81330 65882
rect 81382 65830 81434 65882
rect 81486 65830 81538 65882
rect 111998 65830 112050 65882
rect 112102 65830 112154 65882
rect 112206 65830 112258 65882
rect 1822 65662 1874 65714
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 96638 65046 96690 65098
rect 96742 65046 96794 65098
rect 96846 65046 96898 65098
rect 1822 64430 1874 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 81278 64262 81330 64314
rect 81382 64262 81434 64314
rect 81486 64262 81538 64314
rect 111998 64262 112050 64314
rect 112102 64262 112154 64314
rect 112206 64262 112258 64314
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 96638 63478 96690 63530
rect 96742 63478 96794 63530
rect 96846 63478 96898 63530
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 81278 62694 81330 62746
rect 81382 62694 81434 62746
rect 81486 62694 81538 62746
rect 111998 62694 112050 62746
rect 112102 62694 112154 62746
rect 112206 62694 112258 62746
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 96638 61910 96690 61962
rect 96742 61910 96794 61962
rect 96846 61910 96898 61962
rect 1822 61294 1874 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 81278 61126 81330 61178
rect 81382 61126 81434 61178
rect 81486 61126 81538 61178
rect 111998 61126 112050 61178
rect 112102 61126 112154 61178
rect 112206 61126 112258 61178
rect 118078 60846 118130 60898
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 96638 60342 96690 60394
rect 96742 60342 96794 60394
rect 96846 60342 96898 60394
rect 118078 59838 118130 59890
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 81278 59558 81330 59610
rect 81382 59558 81434 59610
rect 81486 59558 81538 59610
rect 111998 59558 112050 59610
rect 112102 59558 112154 59610
rect 112206 59558 112258 59610
rect 118078 59278 118130 59330
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 96638 58774 96690 58826
rect 96742 58774 96794 58826
rect 96846 58774 96898 58826
rect 1822 58158 1874 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 81278 57990 81330 58042
rect 81382 57990 81434 58042
rect 81486 57990 81538 58042
rect 111998 57990 112050 58042
rect 112102 57990 112154 58042
rect 112206 57990 112258 58042
rect 118078 57710 118130 57762
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 96638 57206 96690 57258
rect 96742 57206 96794 57258
rect 96846 57206 96898 57258
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 81278 56422 81330 56474
rect 81382 56422 81434 56474
rect 81486 56422 81538 56474
rect 111998 56422 112050 56474
rect 112102 56422 112154 56474
rect 112206 56422 112258 56474
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 96638 55638 96690 55690
rect 96742 55638 96794 55690
rect 96846 55638 96898 55690
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 81278 54854 81330 54906
rect 81382 54854 81434 54906
rect 81486 54854 81538 54906
rect 111998 54854 112050 54906
rect 112102 54854 112154 54906
rect 112206 54854 112258 54906
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 96638 54070 96690 54122
rect 96742 54070 96794 54122
rect 96846 54070 96898 54122
rect 118078 53454 118130 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 81278 53286 81330 53338
rect 81382 53286 81434 53338
rect 81486 53286 81538 53338
rect 111998 53286 112050 53338
rect 112102 53286 112154 53338
rect 112206 53286 112258 53338
rect 2158 53118 2210 53170
rect 118078 53006 118130 53058
rect 1822 52894 1874 52946
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 96638 52502 96690 52554
rect 96742 52502 96794 52554
rect 96846 52502 96898 52554
rect 1822 52222 1874 52274
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 81278 51718 81330 51770
rect 81382 51718 81434 51770
rect 81486 51718 81538 51770
rect 111998 51718 112050 51770
rect 112102 51718 112154 51770
rect 112206 51718 112258 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 96638 50934 96690 50986
rect 96742 50934 96794 50986
rect 96846 50934 96898 50986
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 81278 50150 81330 50202
rect 81382 50150 81434 50202
rect 81486 50150 81538 50202
rect 111998 50150 112050 50202
rect 112102 50150 112154 50202
rect 112206 50150 112258 50202
rect 1822 49870 1874 49922
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 96638 49366 96690 49418
rect 96742 49366 96794 49418
rect 96846 49366 96898 49418
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 81278 48582 81330 48634
rect 81382 48582 81434 48634
rect 81486 48582 81538 48634
rect 111998 48582 112050 48634
rect 112102 48582 112154 48634
rect 112206 48582 112258 48634
rect 3054 48190 3106 48242
rect 2046 48078 2098 48130
rect 3502 48078 3554 48130
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 96638 47798 96690 47850
rect 96742 47798 96794 47850
rect 96846 47798 96898 47850
rect 118078 47182 118130 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 81278 47014 81330 47066
rect 81382 47014 81434 47066
rect 81486 47014 81538 47066
rect 111998 47014 112050 47066
rect 112102 47014 112154 47066
rect 112206 47014 112258 47066
rect 1822 46734 1874 46786
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 96638 46230 96690 46282
rect 96742 46230 96794 46282
rect 96846 46230 96898 46282
rect 1934 45838 1986 45890
rect 2158 45614 2210 45666
rect 2606 45614 2658 45666
rect 118078 45614 118130 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 81278 45446 81330 45498
rect 81382 45446 81434 45498
rect 81486 45446 81538 45498
rect 111998 45446 112050 45498
rect 112102 45446 112154 45498
rect 112206 45446 112258 45498
rect 2158 45278 2210 45330
rect 1822 45054 1874 45106
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 96638 44662 96690 44714
rect 96742 44662 96794 44714
rect 96846 44662 96898 44714
rect 1822 44382 1874 44434
rect 118078 44046 118130 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 81278 43878 81330 43930
rect 81382 43878 81434 43930
rect 81486 43878 81538 43930
rect 111998 43878 112050 43930
rect 112102 43878 112154 43930
rect 112206 43878 112258 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 96638 43094 96690 43146
rect 96742 43094 96794 43146
rect 96846 43094 96898 43146
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 81278 42310 81330 42362
rect 81382 42310 81434 42362
rect 81486 42310 81538 42362
rect 111998 42310 112050 42362
rect 112102 42310 112154 42362
rect 112206 42310 112258 42362
rect 1822 42030 1874 42082
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 96638 41526 96690 41578
rect 96742 41526 96794 41578
rect 96846 41526 96898 41578
rect 59950 41022 60002 41074
rect 118078 41022 118130 41074
rect 1822 40910 1874 40962
rect 59390 40910 59442 40962
rect 60286 40910 60338 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 81278 40742 81330 40794
rect 81382 40742 81434 40794
rect 81486 40742 81538 40794
rect 111998 40742 112050 40794
rect 112102 40742 112154 40794
rect 112206 40742 112258 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 96638 39958 96690 40010
rect 96742 39958 96794 40010
rect 96846 39958 96898 40010
rect 1822 39342 1874 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 81278 39174 81330 39226
rect 81382 39174 81434 39226
rect 81486 39174 81538 39226
rect 111998 39174 112050 39226
rect 112102 39174 112154 39226
rect 112206 39174 112258 39226
rect 118078 38894 118130 38946
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 96638 38390 96690 38442
rect 96742 38390 96794 38442
rect 96846 38390 96898 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 81278 37606 81330 37658
rect 81382 37606 81434 37658
rect 81486 37606 81538 37658
rect 111998 37606 112050 37658
rect 112102 37606 112154 37658
rect 112206 37606 112258 37658
rect 1822 37326 1874 37378
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 96638 36822 96690 36874
rect 96742 36822 96794 36874
rect 96846 36822 96898 36874
rect 1822 36206 1874 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 81278 36038 81330 36090
rect 81382 36038 81434 36090
rect 81486 36038 81538 36090
rect 111998 36038 112050 36090
rect 112102 36038 112154 36090
rect 112206 36038 112258 36090
rect 117742 35758 117794 35810
rect 116846 35646 116898 35698
rect 116286 35534 116338 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 96638 35254 96690 35306
rect 96742 35254 96794 35306
rect 96846 35254 96898 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 81278 34470 81330 34522
rect 81382 34470 81434 34522
rect 81486 34470 81538 34522
rect 111998 34470 112050 34522
rect 112102 34470 112154 34522
rect 112206 34470 112258 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 96638 33686 96690 33738
rect 96742 33686 96794 33738
rect 96846 33686 96898 33738
rect 1822 33070 1874 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 81278 32902 81330 32954
rect 81382 32902 81434 32954
rect 81486 32902 81538 32954
rect 111998 32902 112050 32954
rect 112102 32902 112154 32954
rect 112206 32902 112258 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 96638 32118 96690 32170
rect 96742 32118 96794 32170
rect 96846 32118 96898 32170
rect 118078 31502 118130 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 81278 31334 81330 31386
rect 81382 31334 81434 31386
rect 81486 31334 81538 31386
rect 111998 31334 112050 31386
rect 112102 31334 112154 31386
rect 112206 31334 112258 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 96638 30550 96690 30602
rect 96742 30550 96794 30602
rect 96846 30550 96898 30602
rect 1822 29934 1874 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 81278 29766 81330 29818
rect 81382 29766 81434 29818
rect 81486 29766 81538 29818
rect 111998 29766 112050 29818
rect 112102 29766 112154 29818
rect 112206 29766 112258 29818
rect 118078 29486 118130 29538
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 96638 28982 96690 29034
rect 96742 28982 96794 29034
rect 96846 28982 96898 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 81278 28198 81330 28250
rect 81382 28198 81434 28250
rect 81486 28198 81538 28250
rect 111998 28198 112050 28250
rect 112102 28198 112154 28250
rect 112206 28198 112258 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 96638 27414 96690 27466
rect 96742 27414 96794 27466
rect 96846 27414 96898 27466
rect 118078 26798 118130 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 81278 26630 81330 26682
rect 81382 26630 81434 26682
rect 81486 26630 81538 26682
rect 111998 26630 112050 26682
rect 112102 26630 112154 26682
rect 112206 26630 112258 26682
rect 1822 26350 1874 26402
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 96638 25846 96690 25898
rect 96742 25846 96794 25898
rect 96846 25846 96898 25898
rect 118078 25230 118130 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 81278 25062 81330 25114
rect 81382 25062 81434 25114
rect 81486 25062 81538 25114
rect 111998 25062 112050 25114
rect 112102 25062 112154 25114
rect 112206 25062 112258 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 96638 24278 96690 24330
rect 96742 24278 96794 24330
rect 96846 24278 96898 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 81278 23494 81330 23546
rect 81382 23494 81434 23546
rect 81486 23494 81538 23546
rect 111998 23494 112050 23546
rect 112102 23494 112154 23546
rect 112206 23494 112258 23546
rect 1822 23214 1874 23266
rect 118078 23214 118130 23266
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 96638 22710 96690 22762
rect 96742 22710 96794 22762
rect 96846 22710 96898 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 81278 21926 81330 21978
rect 81382 21926 81434 21978
rect 81486 21926 81538 21978
rect 111998 21926 112050 21978
rect 112102 21926 112154 21978
rect 112206 21926 112258 21978
rect 1822 21646 1874 21698
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 96638 21142 96690 21194
rect 96742 21142 96794 21194
rect 96846 21142 96898 21194
rect 118078 20526 118130 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 81278 20358 81330 20410
rect 81382 20358 81434 20410
rect 81486 20358 81538 20410
rect 111998 20358 112050 20410
rect 112102 20358 112154 20410
rect 112206 20358 112258 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 96638 19574 96690 19626
rect 96742 19574 96794 19626
rect 96846 19574 96898 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 81278 18790 81330 18842
rect 81382 18790 81434 18842
rect 81486 18790 81538 18842
rect 111998 18790 112050 18842
rect 112102 18790 112154 18842
rect 112206 18790 112258 18842
rect 1822 18510 1874 18562
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 96638 18006 96690 18058
rect 96742 18006 96794 18058
rect 96846 18006 96898 18058
rect 118078 17502 118130 17554
rect 1822 17390 1874 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 81278 17222 81330 17274
rect 81382 17222 81434 17274
rect 81486 17222 81538 17274
rect 111998 17222 112050 17274
rect 112102 17222 112154 17274
rect 112206 17222 112258 17274
rect 118078 16942 118130 16994
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 96638 16438 96690 16490
rect 96742 16438 96794 16490
rect 96846 16438 96898 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 81278 15654 81330 15706
rect 81382 15654 81434 15706
rect 81486 15654 81538 15706
rect 111998 15654 112050 15706
rect 112102 15654 112154 15706
rect 112206 15654 112258 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 96638 14870 96690 14922
rect 96742 14870 96794 14922
rect 96846 14870 96898 14922
rect 118078 14254 118130 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 81278 14086 81330 14138
rect 81382 14086 81434 14138
rect 81486 14086 81538 14138
rect 111998 14086 112050 14138
rect 112102 14086 112154 14138
rect 112206 14086 112258 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 96638 13302 96690 13354
rect 96742 13302 96794 13354
rect 96846 13302 96898 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 81278 12518 81330 12570
rect 81382 12518 81434 12570
rect 81486 12518 81538 12570
rect 111998 12518 112050 12570
rect 112102 12518 112154 12570
rect 112206 12518 112258 12570
rect 118078 12238 118130 12290
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 96638 11734 96690 11786
rect 96742 11734 96794 11786
rect 96846 11734 96898 11786
rect 1822 11118 1874 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 81278 10950 81330 11002
rect 81382 10950 81434 11002
rect 81486 10950 81538 11002
rect 111998 10950 112050 11002
rect 112102 10950 112154 11002
rect 112206 10950 112258 11002
rect 118078 10670 118130 10722
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 96638 10166 96690 10218
rect 96742 10166 96794 10218
rect 96846 10166 96898 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 81278 9382 81330 9434
rect 81382 9382 81434 9434
rect 81486 9382 81538 9434
rect 111998 9382 112050 9434
rect 112102 9382 112154 9434
rect 112206 9382 112258 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 96638 8598 96690 8650
rect 96742 8598 96794 8650
rect 96846 8598 96898 8650
rect 1822 7982 1874 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 81278 7814 81330 7866
rect 81382 7814 81434 7866
rect 81486 7814 81538 7866
rect 111998 7814 112050 7866
rect 112102 7814 112154 7866
rect 112206 7814 112258 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 96638 7030 96690 7082
rect 96742 7030 96794 7082
rect 96846 7030 96898 7082
rect 1822 6414 1874 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 81278 6246 81330 6298
rect 81382 6246 81434 6298
rect 81486 6246 81538 6298
rect 111998 6246 112050 6298
rect 112102 6246 112154 6298
rect 112206 6246 112258 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 96638 5462 96690 5514
rect 96742 5462 96794 5514
rect 96846 5462 96898 5514
rect 1822 4846 1874 4898
rect 118078 4846 118130 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 81278 4678 81330 4730
rect 81382 4678 81434 4730
rect 81486 4678 81538 4730
rect 111998 4678 112050 4730
rect 112102 4678 112154 4730
rect 112206 4678 112258 4730
rect 1822 4398 1874 4450
rect 117182 4398 117234 4450
rect 118078 4398 118130 4450
rect 116510 4174 116562 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 96638 3894 96690 3946
rect 96742 3894 96794 3946
rect 96846 3894 96898 3946
rect 116846 3502 116898 3554
rect 117742 3390 117794 3442
rect 2270 3278 2322 3330
rect 7646 3278 7698 3330
rect 8318 3278 8370 3330
rect 9662 3278 9714 3330
rect 12350 3278 12402 3330
rect 15038 3278 15090 3330
rect 27134 3278 27186 3330
rect 28366 3278 28418 3330
rect 29822 3278 29874 3330
rect 30494 3278 30546 3330
rect 33182 3278 33234 3330
rect 34526 3278 34578 3330
rect 37214 3278 37266 3330
rect 37886 3278 37938 3330
rect 43262 3278 43314 3330
rect 45278 3278 45330 3330
rect 47966 3278 48018 3330
rect 49310 3278 49362 3330
rect 51886 3278 51938 3330
rect 52782 3278 52834 3330
rect 54014 3278 54066 3330
rect 55358 3278 55410 3330
rect 59390 3278 59442 3330
rect 62750 3278 62802 3330
rect 68462 3278 68514 3330
rect 69134 3278 69186 3330
rect 70142 3278 70194 3330
rect 76302 3278 76354 3330
rect 77534 3278 77586 3330
rect 78878 3278 78930 3330
rect 82910 3278 82962 3330
rect 84926 3278 84978 3330
rect 86270 3278 86322 3330
rect 88062 3278 88114 3330
rect 93662 3278 93714 3330
rect 101054 3278 101106 3330
rect 107662 3278 107714 3330
rect 109790 3278 109842 3330
rect 111582 3278 111634 3330
rect 112478 3278 112530 3330
rect 115838 3278 115890 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 81278 3110 81330 3162
rect 81382 3110 81434 3162
rect 81486 3110 81538 3162
rect 111998 3110 112050 3162
rect 112102 3110 112154 3162
rect 112206 3110 112258 3162
rect 87390 1822 87442 1874
rect 88062 1822 88114 1874
rect 110910 1822 110962 1874
rect 111582 1822 111634 1874
rect 67902 1710 67954 1762
rect 68462 1710 68514 1762
<< metal2 >>
rect 114940 135884 115220 135940
rect 114940 135800 114996 135884
rect 0 135200 112 135800
rect 1344 135200 1456 135800
rect 2688 135200 2800 135800
rect 4032 135200 4144 135800
rect 5376 135200 5488 135800
rect 6720 135200 6832 135800
rect 7392 135200 7504 135800
rect 8736 135200 8848 135800
rect 10080 135200 10192 135800
rect 11424 135200 11536 135800
rect 12768 135200 12880 135800
rect 14112 135200 14224 135800
rect 14784 135200 14896 135800
rect 16128 135200 16240 135800
rect 17472 135200 17584 135800
rect 18816 135200 18928 135800
rect 20160 135200 20272 135800
rect 21504 135200 21616 135800
rect 22176 135200 22288 135800
rect 23520 135200 23632 135800
rect 24864 135200 24976 135800
rect 26208 135200 26320 135800
rect 27552 135200 27664 135800
rect 28896 135200 29008 135800
rect 29568 135200 29680 135800
rect 30912 135200 31024 135800
rect 32256 135200 32368 135800
rect 33600 135200 33712 135800
rect 34944 135200 35056 135800
rect 36288 135200 36400 135800
rect 36960 135200 37072 135800
rect 38304 135200 38416 135800
rect 39648 135200 39760 135800
rect 40992 135200 41104 135800
rect 42336 135200 42448 135800
rect 43680 135200 43792 135800
rect 44352 135200 44464 135800
rect 45696 135200 45808 135800
rect 47040 135200 47152 135800
rect 48384 135200 48496 135800
rect 49728 135200 49840 135800
rect 51072 135200 51184 135800
rect 51744 135200 51856 135800
rect 53088 135200 53200 135800
rect 54432 135200 54544 135800
rect 55776 135200 55888 135800
rect 57120 135200 57232 135800
rect 58464 135200 58576 135800
rect 59808 135200 59920 135800
rect 60480 135200 60592 135800
rect 61824 135200 61936 135800
rect 63168 135200 63280 135800
rect 64512 135200 64624 135800
rect 65856 135200 65968 135800
rect 67200 135200 67312 135800
rect 67872 135200 67984 135800
rect 69216 135200 69328 135800
rect 70560 135200 70672 135800
rect 71904 135200 72016 135800
rect 73248 135200 73360 135800
rect 74592 135200 74704 135800
rect 75264 135200 75376 135800
rect 76608 135200 76720 135800
rect 77952 135200 78064 135800
rect 79296 135200 79408 135800
rect 80640 135200 80752 135800
rect 81984 135200 82096 135800
rect 82656 135200 82768 135800
rect 84000 135200 84112 135800
rect 85344 135200 85456 135800
rect 86688 135200 86800 135800
rect 88032 135200 88144 135800
rect 89376 135200 89488 135800
rect 90048 135200 90160 135800
rect 91392 135200 91504 135800
rect 92736 135200 92848 135800
rect 94080 135200 94192 135800
rect 95424 135200 95536 135800
rect 96768 135200 96880 135800
rect 97440 135200 97552 135800
rect 98784 135200 98896 135800
rect 100128 135200 100240 135800
rect 101472 135200 101584 135800
rect 102816 135200 102928 135800
rect 104160 135200 104272 135800
rect 104832 135200 104944 135800
rect 106176 135200 106288 135800
rect 107520 135200 107632 135800
rect 108864 135200 108976 135800
rect 110208 135200 110320 135800
rect 111552 135200 111664 135800
rect 112224 135200 112336 135800
rect 113568 135200 113680 135800
rect 114912 135200 115024 135800
rect 115164 135492 115220 135884
rect 115164 135436 115556 135492
rect 2492 134484 2548 134494
rect 1820 133140 1876 133150
rect 1820 132018 1876 133084
rect 1820 131966 1822 132018
rect 1874 131966 1876 132018
rect 1820 131954 1876 131966
rect 2492 132018 2548 134428
rect 4476 132524 4740 132534
rect 4532 132468 4580 132524
rect 4636 132468 4684 132524
rect 4476 132458 4740 132468
rect 2492 131966 2494 132018
rect 2546 131966 2548 132018
rect 2492 131954 2548 131966
rect 10108 132020 10164 135200
rect 10332 132020 10388 132030
rect 10108 132018 10388 132020
rect 10108 131966 10334 132018
rect 10386 131966 10388 132018
rect 10108 131964 10388 131966
rect 11452 132020 11508 135200
rect 11676 132020 11732 132030
rect 11452 132018 11732 132020
rect 11452 131966 11678 132018
rect 11730 131966 11732 132018
rect 11452 131964 11732 131966
rect 10332 131954 10388 131964
rect 11676 131954 11732 131964
rect 12796 132020 12852 135200
rect 20188 132244 20244 135200
rect 20188 132178 20244 132188
rect 22092 132244 22148 132254
rect 22092 132150 22148 132188
rect 21420 132130 21476 132142
rect 21420 132078 21422 132130
rect 21474 132078 21476 132130
rect 12796 131954 12852 131964
rect 13580 132020 13636 132030
rect 13580 131926 13636 131964
rect 20636 131908 20692 131918
rect 21420 131908 21476 132078
rect 23548 132020 23604 135200
rect 23772 132020 23828 132030
rect 23548 132018 23828 132020
rect 23548 131966 23774 132018
rect 23826 131966 23828 132018
rect 23548 131964 23828 131966
rect 26236 132020 26292 135200
rect 26460 132020 26516 132030
rect 26236 132018 26516 132020
rect 26236 131966 26462 132018
rect 26514 131966 26516 132018
rect 26236 131964 26516 131966
rect 27580 132020 27636 135200
rect 27804 132020 27860 132030
rect 27580 132018 27860 132020
rect 27580 131966 27806 132018
rect 27858 131966 27860 132018
rect 27580 131964 27860 131966
rect 29596 132020 29652 135200
rect 29820 132020 29876 132030
rect 29596 132018 29876 132020
rect 29596 131966 29822 132018
rect 29874 131966 29876 132018
rect 29596 131964 29876 131966
rect 30940 132020 30996 135200
rect 35196 132524 35460 132534
rect 35252 132468 35300 132524
rect 35356 132468 35404 132524
rect 35196 132458 35460 132468
rect 31164 132020 31220 132030
rect 30940 132018 31220 132020
rect 30940 131966 31166 132018
rect 31218 131966 31220 132018
rect 30940 131964 31220 131966
rect 23772 131954 23828 131964
rect 26460 131954 26516 131964
rect 27804 131954 27860 131964
rect 29820 131954 29876 131964
rect 31164 131954 31220 131964
rect 36316 132018 36372 135200
rect 36316 131966 36318 132018
rect 36370 131966 36372 132018
rect 36316 131954 36372 131966
rect 36988 132020 37044 135200
rect 37212 132020 37268 132030
rect 36988 132018 37268 132020
rect 36988 131966 37214 132018
rect 37266 131966 37268 132018
rect 36988 131964 37268 131966
rect 39676 132020 39732 135200
rect 39900 132020 39956 132030
rect 39676 132018 39956 132020
rect 39676 131966 39902 132018
rect 39954 131966 39956 132018
rect 39676 131964 39956 131966
rect 45724 132020 45780 135200
rect 45948 132020 46004 132030
rect 45724 132018 46004 132020
rect 45724 131966 45950 132018
rect 46002 131966 46004 132018
rect 45724 131964 46004 131966
rect 51100 132020 51156 135200
rect 51324 132020 51380 132030
rect 51100 132018 51380 132020
rect 51100 131966 51326 132018
rect 51378 131966 51380 132018
rect 51100 131964 51380 131966
rect 53116 132020 53172 135200
rect 53340 132020 53396 132030
rect 53116 132018 53396 132020
rect 53116 131966 53342 132018
rect 53394 131966 53396 132018
rect 53116 131964 53396 131966
rect 54460 132020 54516 135200
rect 54684 132020 54740 132030
rect 54460 132018 54740 132020
rect 54460 131966 54686 132018
rect 54738 131966 54740 132018
rect 54460 131964 54740 131966
rect 58492 132020 58548 135200
rect 59836 132242 59892 135200
rect 60508 132690 60564 135200
rect 60508 132638 60510 132690
rect 60562 132638 60564 132690
rect 60508 132626 60564 132638
rect 61516 132690 61572 132702
rect 61516 132638 61518 132690
rect 61570 132638 61572 132690
rect 59836 132190 59838 132242
rect 59890 132190 59892 132242
rect 59836 132132 59892 132190
rect 59836 132066 59892 132076
rect 60844 132132 60900 132142
rect 60844 132038 60900 132076
rect 58716 132020 58772 132030
rect 58492 132018 58772 132020
rect 58492 131966 58718 132018
rect 58770 131966 58772 132018
rect 58492 131964 58772 131966
rect 37212 131954 37268 131964
rect 39900 131954 39956 131964
rect 45948 131954 46004 131964
rect 51324 131954 51380 131964
rect 53340 131954 53396 131964
rect 54684 131954 54740 131964
rect 58716 131954 58772 131964
rect 61516 132018 61572 132638
rect 61516 131966 61518 132018
rect 61570 131966 61572 132018
rect 61516 131954 61572 131966
rect 63196 132020 63252 135200
rect 63420 132020 63476 132030
rect 63196 132018 63476 132020
rect 63196 131966 63422 132018
rect 63474 131966 63476 132018
rect 63196 131964 63476 131966
rect 64540 132020 64596 135200
rect 65884 133700 65940 135200
rect 65772 133644 65940 133700
rect 65772 132356 65828 133644
rect 65916 132524 66180 132534
rect 65972 132468 66020 132524
rect 66076 132468 66124 132524
rect 65916 132458 66180 132468
rect 65772 132300 66164 132356
rect 64764 132020 64820 132030
rect 64540 132018 64820 132020
rect 64540 131966 64766 132018
rect 64818 131966 64820 132018
rect 64540 131964 64820 131966
rect 63420 131954 63476 131964
rect 64764 131954 64820 131964
rect 66108 132018 66164 132300
rect 66108 131966 66110 132018
rect 66162 131966 66164 132018
rect 66108 131954 66164 131966
rect 67228 132020 67284 135200
rect 67452 132020 67508 132030
rect 67228 132018 67508 132020
rect 67228 131966 67454 132018
rect 67506 131966 67508 132018
rect 67228 131964 67508 131966
rect 69244 132020 69300 135200
rect 69468 132020 69524 132030
rect 69244 132018 69524 132020
rect 69244 131966 69470 132018
rect 69522 131966 69524 132018
rect 69244 131964 69524 131966
rect 67452 131954 67508 131964
rect 69468 131954 69524 131964
rect 71932 132020 71988 135200
rect 71932 131954 71988 131964
rect 72380 132020 72436 132030
rect 73276 132020 73332 135200
rect 73500 132020 73556 132030
rect 73276 132018 73556 132020
rect 73276 131966 73502 132018
rect 73554 131966 73556 132018
rect 73276 131964 73556 131966
rect 74620 132020 74676 135200
rect 74844 132020 74900 132030
rect 74620 132018 74900 132020
rect 74620 131966 74846 132018
rect 74898 131966 74900 132018
rect 74620 131964 74900 131966
rect 72380 131926 72436 131964
rect 73500 131954 73556 131964
rect 74844 131954 74900 131964
rect 75292 132020 75348 135200
rect 75292 131954 75348 131964
rect 76300 132020 76356 132030
rect 80668 132020 80724 135200
rect 80892 132020 80948 132030
rect 80668 132018 80948 132020
rect 80668 131966 80894 132018
rect 80946 131966 80948 132018
rect 80668 131964 80948 131966
rect 82012 132020 82068 135200
rect 82236 132020 82292 132030
rect 82012 132018 82292 132020
rect 82012 131966 82238 132018
rect 82290 131966 82292 132018
rect 82012 131964 82292 131966
rect 84028 132020 84084 135200
rect 84252 132020 84308 132030
rect 84028 132018 84308 132020
rect 84028 131966 84254 132018
rect 84306 131966 84308 132018
rect 84028 131964 84308 131966
rect 85372 132020 85428 135200
rect 85596 132020 85652 132030
rect 85372 132018 85652 132020
rect 85372 131966 85598 132018
rect 85650 131966 85652 132018
rect 85372 131964 85652 131966
rect 88060 132020 88116 135200
rect 88284 132020 88340 132030
rect 88060 132018 88340 132020
rect 88060 131966 88286 132018
rect 88338 131966 88340 132018
rect 88060 131964 88340 131966
rect 89404 132020 89460 135200
rect 89628 132020 89684 132030
rect 89404 132018 89684 132020
rect 89404 131966 89630 132018
rect 89682 131966 89684 132018
rect 89404 131964 89684 131966
rect 76300 131926 76356 131964
rect 80892 131954 80948 131964
rect 82236 131954 82292 131964
rect 84252 131954 84308 131964
rect 85596 131954 85652 131964
rect 88284 131954 88340 131964
rect 89628 131954 89684 131964
rect 95452 132020 95508 135200
rect 102844 132690 102900 135200
rect 102844 132638 102846 132690
rect 102898 132638 102900 132690
rect 102844 132626 102900 132638
rect 103740 132690 103796 132702
rect 103740 132638 103742 132690
rect 103794 132638 103796 132690
rect 96636 132524 96900 132534
rect 96692 132468 96740 132524
rect 96796 132468 96844 132524
rect 96636 132458 96900 132468
rect 95452 131954 95508 131964
rect 95900 132020 95956 132030
rect 95900 131926 95956 131964
rect 103740 132018 103796 132638
rect 103740 131966 103742 132018
rect 103794 131966 103796 132018
rect 103740 131954 103796 131966
rect 104188 132020 104244 135200
rect 104412 132020 104468 132030
rect 104188 132018 104468 132020
rect 104188 131966 104414 132018
rect 104466 131966 104468 132018
rect 104188 131964 104468 131966
rect 108892 132020 108948 135200
rect 109116 132020 109172 132030
rect 108892 132018 109172 132020
rect 108892 131966 109118 132018
rect 109170 131966 109172 132018
rect 108892 131964 109172 131966
rect 104412 131954 104468 131964
rect 109116 131954 109172 131964
rect 115500 132018 115556 135436
rect 116256 135200 116368 135800
rect 117600 135200 117712 135800
rect 118944 135200 119056 135800
rect 119616 135200 119728 135800
rect 115500 131966 115502 132018
rect 115554 131966 115556 132018
rect 115500 131954 115556 131966
rect 116284 132020 116340 135200
rect 117292 132468 117348 132478
rect 116508 132020 116564 132030
rect 116284 132018 116564 132020
rect 116284 131966 116510 132018
rect 116562 131966 116564 132018
rect 116284 131964 116564 131966
rect 116508 131954 116564 131964
rect 117292 132018 117348 132412
rect 117292 131966 117294 132018
rect 117346 131966 117348 132018
rect 117292 131954 117348 131966
rect 117628 132020 117684 135200
rect 117852 132020 117908 132030
rect 117628 132018 117908 132020
rect 117628 131966 117854 132018
rect 117906 131966 117908 132018
rect 117628 131964 117908 131966
rect 117852 131954 117908 131964
rect 20636 131906 21476 131908
rect 20636 131854 20638 131906
rect 20690 131854 21476 131906
rect 20636 131852 21476 131854
rect 20636 131842 20692 131852
rect 19836 131740 20100 131750
rect 19892 131684 19940 131740
rect 19996 131684 20044 131740
rect 19836 131674 20100 131684
rect 4476 130956 4740 130966
rect 4532 130900 4580 130956
rect 4636 130900 4684 130956
rect 4476 130890 4740 130900
rect 1820 130452 1876 130462
rect 1820 130358 1876 130396
rect 19836 130172 20100 130182
rect 19892 130116 19940 130172
rect 19996 130116 20044 130172
rect 19836 130106 20100 130116
rect 4476 129388 4740 129398
rect 4532 129332 4580 129388
rect 4636 129332 4684 129388
rect 4476 129322 4740 129332
rect 19836 128604 20100 128614
rect 19892 128548 19940 128604
rect 19996 128548 20044 128604
rect 19836 128538 20100 128548
rect 1820 128322 1876 128334
rect 1820 128270 1822 128322
rect 1874 128270 1876 128322
rect 1820 127764 1876 128270
rect 4476 127820 4740 127830
rect 4532 127764 4580 127820
rect 4636 127764 4684 127820
rect 4476 127754 4740 127764
rect 1820 127698 1876 127708
rect 1820 127202 1876 127214
rect 1820 127150 1822 127202
rect 1874 127150 1876 127202
rect 1820 127092 1876 127150
rect 1820 127026 1876 127036
rect 19836 127036 20100 127046
rect 19892 126980 19940 127036
rect 19996 126980 20044 127036
rect 19836 126970 20100 126980
rect 4476 126252 4740 126262
rect 4532 126196 4580 126252
rect 4636 126196 4684 126252
rect 4476 126186 4740 126196
rect 19836 125468 20100 125478
rect 19892 125412 19940 125468
rect 19996 125412 20044 125468
rect 19836 125402 20100 125412
rect 1820 125186 1876 125198
rect 1820 125134 1822 125186
rect 1874 125134 1876 125186
rect 1820 124404 1876 125134
rect 4476 124684 4740 124694
rect 4532 124628 4580 124684
rect 4636 124628 4684 124684
rect 4476 124618 4740 124628
rect 1820 124338 1876 124348
rect 19836 123900 20100 123910
rect 19892 123844 19940 123900
rect 19996 123844 20044 123900
rect 19836 123834 20100 123844
rect 1820 123618 1876 123630
rect 1820 123566 1822 123618
rect 1874 123566 1876 123618
rect 1820 123060 1876 123566
rect 4476 123116 4740 123126
rect 4532 123060 4580 123116
rect 4636 123060 4684 123116
rect 4476 123050 4740 123060
rect 1820 122994 1876 123004
rect 19836 122332 20100 122342
rect 19892 122276 19940 122332
rect 19996 122276 20044 122332
rect 19836 122266 20100 122276
rect 1820 122050 1876 122062
rect 1820 121998 1822 122050
rect 1874 121998 1876 122050
rect 1820 121716 1876 121998
rect 1820 121650 1876 121660
rect 4476 121548 4740 121558
rect 4532 121492 4580 121548
rect 4636 121492 4684 121548
rect 4476 121482 4740 121492
rect 19836 120764 20100 120774
rect 19892 120708 19940 120764
rect 19996 120708 20044 120764
rect 19836 120698 20100 120708
rect 4476 119980 4740 119990
rect 4532 119924 4580 119980
rect 4636 119924 4684 119980
rect 4476 119914 4740 119924
rect 19836 119196 20100 119206
rect 19892 119140 19940 119196
rect 19996 119140 20044 119196
rect 19836 119130 20100 119140
rect 4476 118412 4740 118422
rect 4532 118356 4580 118412
rect 4636 118356 4684 118412
rect 4476 118346 4740 118356
rect 19836 117628 20100 117638
rect 19892 117572 19940 117628
rect 19996 117572 20044 117628
rect 19836 117562 20100 117572
rect 1820 117346 1876 117358
rect 1820 117294 1822 117346
rect 1874 117294 1876 117346
rect 1820 117012 1876 117294
rect 1820 116946 1876 116956
rect 4476 116844 4740 116854
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4476 116778 4740 116788
rect 19836 116060 20100 116070
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 19836 115994 20100 116004
rect 4476 115276 4740 115286
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4476 115210 4740 115220
rect 19836 114492 20100 114502
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 19836 114426 20100 114436
rect 4476 113708 4740 113718
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4476 113642 4740 113652
rect 19836 112924 20100 112934
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 19836 112858 20100 112868
rect 4476 112140 4740 112150
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4476 112074 4740 112084
rect 1820 111522 1876 111534
rect 1820 111470 1822 111522
rect 1874 111470 1876 111522
rect 1820 110964 1876 111470
rect 19836 111356 20100 111366
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 19836 111290 20100 111300
rect 1820 110898 1876 110908
rect 4476 110572 4740 110582
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4476 110506 4740 110516
rect 1820 109954 1876 109966
rect 1820 109902 1822 109954
rect 1874 109902 1876 109954
rect 1820 109620 1876 109902
rect 19836 109788 20100 109798
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 19836 109722 20100 109732
rect 1820 109554 1876 109564
rect 4476 109004 4740 109014
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4476 108938 4740 108948
rect 19836 108220 20100 108230
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 19836 108154 20100 108164
rect 4476 107436 4740 107446
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4476 107370 4740 107380
rect 19836 106652 20100 106662
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 19836 106586 20100 106596
rect 4476 105868 4740 105878
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4476 105802 4740 105812
rect 1820 105250 1876 105262
rect 1820 105198 1822 105250
rect 1874 105198 1876 105250
rect 1820 104916 1876 105198
rect 19836 105084 20100 105094
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 19836 105018 20100 105028
rect 1820 104850 1876 104860
rect 4476 104300 4740 104310
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4476 104234 4740 104244
rect 19836 103516 20100 103526
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 19836 103450 20100 103460
rect 4476 102732 4740 102742
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4476 102666 4740 102676
rect 19836 101948 20100 101958
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 19836 101882 20100 101892
rect 1820 101666 1876 101678
rect 1820 101614 1822 101666
rect 1874 101614 1876 101666
rect 1820 100884 1876 101614
rect 4476 101164 4740 101174
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4476 101098 4740 101108
rect 1820 100818 1876 100828
rect 19836 100380 20100 100390
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 19836 100314 20100 100324
rect 4476 99596 4740 99606
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4476 99530 4740 99540
rect 19836 98812 20100 98822
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 19836 98746 20100 98756
rect 4476 98028 4740 98038
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4476 97962 4740 97972
rect 19836 97244 20100 97254
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 19836 97178 20100 97188
rect 1820 96962 1876 96974
rect 1820 96910 1822 96962
rect 1874 96910 1876 96962
rect 1820 96180 1876 96910
rect 4476 96460 4740 96470
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4476 96394 4740 96404
rect 1820 96114 1876 96124
rect 19836 95676 20100 95686
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 19836 95610 20100 95620
rect 1820 95394 1876 95406
rect 1820 95342 1822 95394
rect 1874 95342 1876 95394
rect 1820 94836 1876 95342
rect 4476 94892 4740 94902
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4476 94826 4740 94836
rect 1820 94770 1876 94780
rect 19836 94108 20100 94118
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 19836 94042 20100 94052
rect 4476 93324 4740 93334
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4476 93258 4740 93268
rect 1820 92706 1876 92718
rect 1820 92654 1822 92706
rect 1874 92654 1876 92706
rect 1820 92148 1876 92654
rect 19836 92540 20100 92550
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 19836 92474 20100 92484
rect 1820 92082 1876 92092
rect 4476 91756 4740 91766
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4476 91690 4740 91700
rect 1820 91138 1876 91150
rect 1820 91086 1822 91138
rect 1874 91086 1876 91138
rect 1820 90804 1876 91086
rect 19836 90972 20100 90982
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 19836 90906 20100 90916
rect 1820 90738 1876 90748
rect 2156 90692 2212 90702
rect 1932 90690 2212 90692
rect 1932 90638 2158 90690
rect 2210 90638 2212 90690
rect 1932 90636 2212 90638
rect 1820 90578 1876 90590
rect 1820 90526 1822 90578
rect 1874 90526 1876 90578
rect 1820 90132 1876 90526
rect 1820 89906 1876 90076
rect 1820 89854 1822 89906
rect 1874 89854 1876 89906
rect 1820 89842 1876 89854
rect 1820 83298 1876 83310
rect 1820 83246 1822 83298
rect 1874 83246 1876 83298
rect 1820 82740 1876 83246
rect 1820 82674 1876 82684
rect 1820 78034 1876 78046
rect 1820 77982 1822 78034
rect 1874 77982 1876 78034
rect 1820 77364 1876 77982
rect 1820 77270 1876 77308
rect 1820 73442 1876 73454
rect 1820 73390 1822 73442
rect 1874 73390 1876 73442
rect 1820 72660 1876 73390
rect 1820 72594 1876 72604
rect 1932 67172 1988 90636
rect 2156 90626 2212 90636
rect 4476 90188 4740 90198
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4476 90122 4740 90132
rect 19836 89404 20100 89414
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 19836 89338 20100 89348
rect 4476 88620 4740 88630
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4476 88554 4740 88564
rect 19836 87836 20100 87846
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 19836 87770 20100 87780
rect 4476 87052 4740 87062
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4476 86986 4740 86996
rect 19836 86268 20100 86278
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 19836 86202 20100 86212
rect 4476 85484 4740 85494
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4476 85418 4740 85428
rect 2828 85090 2884 85102
rect 2828 85038 2830 85090
rect 2882 85038 2884 85090
rect 2156 84978 2212 84990
rect 2156 84926 2158 84978
rect 2210 84926 2212 84978
rect 2156 84756 2212 84926
rect 2156 84690 2212 84700
rect 2828 84868 2884 85038
rect 2492 83412 2548 83422
rect 2492 83318 2548 83356
rect 2156 78148 2212 78158
rect 2156 78146 2660 78148
rect 2156 78094 2158 78146
rect 2210 78094 2660 78146
rect 2156 78092 2660 78094
rect 2156 78082 2212 78092
rect 2604 68852 2660 78092
rect 2604 68738 2660 68796
rect 2604 68686 2606 68738
rect 2658 68686 2660 68738
rect 2604 68674 2660 68686
rect 2716 68402 2772 68414
rect 2716 68350 2718 68402
rect 2770 68350 2772 68402
rect 1932 67058 1988 67116
rect 1932 67006 1934 67058
rect 1986 67006 1988 67058
rect 1932 66994 1988 67006
rect 2044 67732 2100 67742
rect 2492 67732 2548 67742
rect 2044 67730 2548 67732
rect 2044 67678 2046 67730
rect 2098 67678 2494 67730
rect 2546 67678 2548 67730
rect 2044 67676 2548 67678
rect 1820 66612 1876 66622
rect 1820 66274 1876 66556
rect 1820 66222 1822 66274
rect 1874 66222 1876 66274
rect 1820 65714 1876 66222
rect 1820 65662 1822 65714
rect 1874 65662 1876 65714
rect 1820 65650 1876 65662
rect 1820 64482 1876 64494
rect 1820 64430 1822 64482
rect 1874 64430 1876 64482
rect 1820 63924 1876 64430
rect 1820 63858 1876 63868
rect 1820 61346 1876 61358
rect 1820 61294 1822 61346
rect 1874 61294 1876 61346
rect 1820 61236 1876 61294
rect 1820 61170 1876 61180
rect 1820 58210 1876 58222
rect 1820 58158 1822 58210
rect 1874 58158 1876 58210
rect 1820 57876 1876 58158
rect 1820 57810 1876 57820
rect 2044 55468 2100 67676
rect 2492 67666 2548 67676
rect 2716 67620 2772 68350
rect 2828 67730 2884 84812
rect 3500 84868 3556 84878
rect 3500 84774 3556 84812
rect 19836 84700 20100 84710
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 19836 84634 20100 84644
rect 4476 83916 4740 83926
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4476 83850 4740 83860
rect 19836 83132 20100 83142
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 19836 83066 20100 83076
rect 4476 82348 4740 82358
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4476 82282 4740 82292
rect 19836 81564 20100 81574
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 19836 81498 20100 81508
rect 4476 80780 4740 80790
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4476 80714 4740 80724
rect 19836 79996 20100 80006
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 19836 79930 20100 79940
rect 4476 79212 4740 79222
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4476 79146 4740 79156
rect 19836 78428 20100 78438
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 19836 78362 20100 78372
rect 4476 77644 4740 77654
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4476 77578 4740 77588
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 3164 68852 3220 68862
rect 3164 68758 3220 68796
rect 20076 68852 20132 68862
rect 20076 68758 20132 68796
rect 21420 68852 21476 131852
rect 60620 131906 60676 131918
rect 60620 131854 60622 131906
rect 60674 131854 60676 131906
rect 50556 131740 50820 131750
rect 50612 131684 50660 131740
rect 50716 131684 50764 131740
rect 50556 131674 50820 131684
rect 35196 130956 35460 130966
rect 35252 130900 35300 130956
rect 35356 130900 35404 130956
rect 35196 130890 35460 130900
rect 50556 130172 50820 130182
rect 50612 130116 50660 130172
rect 50716 130116 50764 130172
rect 50556 130106 50820 130116
rect 35196 129388 35460 129398
rect 35252 129332 35300 129388
rect 35356 129332 35404 129388
rect 35196 129322 35460 129332
rect 50556 128604 50820 128614
rect 50612 128548 50660 128604
rect 50716 128548 50764 128604
rect 50556 128538 50820 128548
rect 35196 127820 35460 127830
rect 35252 127764 35300 127820
rect 35356 127764 35404 127820
rect 35196 127754 35460 127764
rect 50556 127036 50820 127046
rect 50612 126980 50660 127036
rect 50716 126980 50764 127036
rect 50556 126970 50820 126980
rect 35196 126252 35460 126262
rect 35252 126196 35300 126252
rect 35356 126196 35404 126252
rect 35196 126186 35460 126196
rect 50556 125468 50820 125478
rect 50612 125412 50660 125468
rect 50716 125412 50764 125468
rect 50556 125402 50820 125412
rect 35196 124684 35460 124694
rect 35252 124628 35300 124684
rect 35356 124628 35404 124684
rect 35196 124618 35460 124628
rect 50556 123900 50820 123910
rect 50612 123844 50660 123900
rect 50716 123844 50764 123900
rect 50556 123834 50820 123844
rect 35196 123116 35460 123126
rect 35252 123060 35300 123116
rect 35356 123060 35404 123116
rect 35196 123050 35460 123060
rect 50556 122332 50820 122342
rect 50612 122276 50660 122332
rect 50716 122276 50764 122332
rect 50556 122266 50820 122276
rect 35196 121548 35460 121558
rect 35252 121492 35300 121548
rect 35356 121492 35404 121548
rect 35196 121482 35460 121492
rect 50556 120764 50820 120774
rect 50612 120708 50660 120764
rect 50716 120708 50764 120764
rect 50556 120698 50820 120708
rect 35196 119980 35460 119990
rect 35252 119924 35300 119980
rect 35356 119924 35404 119980
rect 35196 119914 35460 119924
rect 50556 119196 50820 119206
rect 50612 119140 50660 119196
rect 50716 119140 50764 119196
rect 50556 119130 50820 119140
rect 35196 118412 35460 118422
rect 35252 118356 35300 118412
rect 35356 118356 35404 118412
rect 35196 118346 35460 118356
rect 50556 117628 50820 117638
rect 50612 117572 50660 117628
rect 50716 117572 50764 117628
rect 50556 117562 50820 117572
rect 35196 116844 35460 116854
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35196 116778 35460 116788
rect 50556 116060 50820 116070
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50556 115994 50820 116004
rect 35196 115276 35460 115286
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35196 115210 35460 115220
rect 50556 114492 50820 114502
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50556 114426 50820 114436
rect 35196 113708 35460 113718
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35196 113642 35460 113652
rect 50556 112924 50820 112934
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50556 112858 50820 112868
rect 35196 112140 35460 112150
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35196 112074 35460 112084
rect 50556 111356 50820 111366
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50556 111290 50820 111300
rect 35196 110572 35460 110582
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35196 110506 35460 110516
rect 50556 109788 50820 109798
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50556 109722 50820 109732
rect 35196 109004 35460 109014
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35196 108938 35460 108948
rect 50556 108220 50820 108230
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50556 108154 50820 108164
rect 35196 107436 35460 107446
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35196 107370 35460 107380
rect 50556 106652 50820 106662
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50556 106586 50820 106596
rect 35196 105868 35460 105878
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35196 105802 35460 105812
rect 50556 105084 50820 105094
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50556 105018 50820 105028
rect 35196 104300 35460 104310
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35196 104234 35460 104244
rect 50556 103516 50820 103526
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50556 103450 50820 103460
rect 35196 102732 35460 102742
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35196 102666 35460 102676
rect 50556 101948 50820 101958
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50556 101882 50820 101892
rect 35196 101164 35460 101174
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35196 101098 35460 101108
rect 50556 100380 50820 100390
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50556 100314 50820 100324
rect 35196 99596 35460 99606
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35196 99530 35460 99540
rect 50556 98812 50820 98822
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50556 98746 50820 98756
rect 35196 98028 35460 98038
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35196 97962 35460 97972
rect 50556 97244 50820 97254
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50556 97178 50820 97188
rect 35196 96460 35460 96470
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35196 96394 35460 96404
rect 50556 95676 50820 95686
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50556 95610 50820 95620
rect 35196 94892 35460 94902
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35196 94826 35460 94836
rect 50556 94108 50820 94118
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50556 94042 50820 94052
rect 35196 93324 35460 93334
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35196 93258 35460 93268
rect 50556 92540 50820 92550
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50556 92474 50820 92484
rect 35196 91756 35460 91766
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35196 91690 35460 91700
rect 50556 90972 50820 90982
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50556 90906 50820 90916
rect 35196 90188 35460 90198
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35196 90122 35460 90132
rect 50556 89404 50820 89414
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50556 89338 50820 89348
rect 35196 88620 35460 88630
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35196 88554 35460 88564
rect 50556 87836 50820 87846
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50556 87770 50820 87780
rect 35196 87052 35460 87062
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35196 86986 35460 86996
rect 50556 86268 50820 86278
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50556 86202 50820 86212
rect 35196 85484 35460 85494
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35196 85418 35460 85428
rect 50556 84700 50820 84710
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50556 84634 50820 84644
rect 35196 83916 35460 83926
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35196 83850 35460 83860
rect 50556 83132 50820 83142
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50556 83066 50820 83076
rect 35196 82348 35460 82358
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35196 82282 35460 82292
rect 50556 81564 50820 81574
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50556 81498 50820 81508
rect 35196 80780 35460 80790
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35196 80714 35460 80724
rect 50556 79996 50820 80006
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50556 79930 50820 79940
rect 35196 79212 35460 79222
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35196 79146 35460 79156
rect 50556 78428 50820 78438
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50556 78362 50820 78372
rect 35196 77644 35460 77654
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35196 77578 35460 77588
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 21420 68786 21476 68796
rect 19964 68516 20020 68526
rect 19964 68422 20020 68460
rect 20636 68516 20692 68526
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 3388 67844 3444 67854
rect 4060 67844 4116 67854
rect 3388 67842 4116 67844
rect 3388 67790 3390 67842
rect 3442 67790 4062 67842
rect 4114 67790 4116 67842
rect 3388 67788 4116 67790
rect 3388 67778 3444 67788
rect 2828 67678 2830 67730
rect 2882 67678 2884 67730
rect 2828 67666 2884 67678
rect 2716 67554 2772 67564
rect 3500 67620 3556 67630
rect 3500 67526 3556 67564
rect 3724 67618 3780 67630
rect 3724 67566 3726 67618
rect 3778 67566 3780 67618
rect 2268 67058 2324 67070
rect 2268 67006 2270 67058
rect 2322 67006 2324 67058
rect 2156 66164 2212 66174
rect 2268 66164 2324 67006
rect 3724 67060 3780 67566
rect 3724 66994 3780 67004
rect 2156 66162 2324 66164
rect 2156 66110 2158 66162
rect 2210 66110 2324 66162
rect 2156 66108 2324 66110
rect 2156 66098 2212 66108
rect 2044 55412 2212 55468
rect 2156 53170 2212 55412
rect 2156 53118 2158 53170
rect 2210 53118 2212 53170
rect 2156 53106 2212 53118
rect 1820 52946 1876 52958
rect 1820 52894 1822 52946
rect 1874 52894 1876 52946
rect 1820 52500 1876 52894
rect 1820 52274 1876 52444
rect 1820 52222 1822 52274
rect 1874 52222 1876 52274
rect 1820 52210 1876 52222
rect 1820 49922 1876 49934
rect 1820 49870 1822 49922
rect 1874 49870 1876 49922
rect 1820 49140 1876 49870
rect 1820 49074 1876 49084
rect 3052 48242 3108 48254
rect 3052 48190 3054 48242
rect 3106 48190 3108 48242
rect 2044 48130 2100 48142
rect 2044 48078 2046 48130
rect 2098 48078 2100 48130
rect 2044 47796 2100 48078
rect 3052 48132 3108 48190
rect 3052 48066 3108 48076
rect 3500 48132 3556 48142
rect 3500 48038 3556 48076
rect 2044 47730 2100 47740
rect 1820 46786 1876 46798
rect 1820 46734 1822 46786
rect 1874 46734 1876 46786
rect 1820 46452 1876 46734
rect 1820 46386 1876 46396
rect 1932 45890 1988 45902
rect 1932 45838 1934 45890
rect 1986 45838 1988 45890
rect 1820 45106 1876 45118
rect 1820 45054 1822 45106
rect 1874 45054 1876 45106
rect 1820 44436 1876 45054
rect 1932 45108 1988 45838
rect 2156 45668 2212 45678
rect 2156 45666 2324 45668
rect 2156 45614 2158 45666
rect 2210 45614 2324 45666
rect 2156 45612 2324 45614
rect 2156 45602 2212 45612
rect 2156 45332 2212 45342
rect 2156 45238 2212 45276
rect 1932 45042 1988 45052
rect 1820 44342 1876 44380
rect 1820 42082 1876 42094
rect 1820 42030 1822 42082
rect 1874 42030 1876 42082
rect 1820 41748 1876 42030
rect 1820 41682 1876 41692
rect 1820 40962 1876 40974
rect 1820 40910 1822 40962
rect 1874 40910 1876 40962
rect 1820 40404 1876 40910
rect 2268 40964 2324 45612
rect 2604 45666 2660 45678
rect 2604 45614 2606 45666
rect 2658 45614 2660 45666
rect 2604 45108 2660 45614
rect 4060 45332 4116 67788
rect 5068 67620 5124 67630
rect 4620 67060 4676 67070
rect 4620 66966 4676 67004
rect 5068 67058 5124 67564
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 6300 67172 6356 67182
rect 6300 67078 6356 67116
rect 5068 67006 5070 67058
rect 5122 67006 5124 67058
rect 5068 66994 5124 67006
rect 5852 66836 5908 66846
rect 5852 66742 5908 66780
rect 20636 66836 20692 68460
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 59612 67956 59668 67966
rect 59612 67842 59668 67900
rect 60060 67956 60116 67966
rect 60060 67862 60116 67900
rect 60620 67956 60676 131854
rect 81276 131740 81540 131750
rect 81332 131684 81380 131740
rect 81436 131684 81484 131740
rect 81276 131674 81540 131684
rect 111996 131740 112260 131750
rect 112052 131684 112100 131740
rect 112156 131684 112204 131740
rect 111996 131674 112260 131684
rect 65916 130956 66180 130966
rect 65972 130900 66020 130956
rect 66076 130900 66124 130956
rect 65916 130890 66180 130900
rect 96636 130956 96900 130966
rect 96692 130900 96740 130956
rect 96796 130900 96844 130956
rect 96636 130890 96900 130900
rect 81276 130172 81540 130182
rect 81332 130116 81380 130172
rect 81436 130116 81484 130172
rect 81276 130106 81540 130116
rect 111996 130172 112260 130182
rect 112052 130116 112100 130172
rect 112156 130116 112204 130172
rect 111996 130106 112260 130116
rect 65916 129388 66180 129398
rect 65972 129332 66020 129388
rect 66076 129332 66124 129388
rect 65916 129322 66180 129332
rect 96636 129388 96900 129398
rect 96692 129332 96740 129388
rect 96796 129332 96844 129388
rect 96636 129322 96900 129332
rect 81276 128604 81540 128614
rect 81332 128548 81380 128604
rect 81436 128548 81484 128604
rect 81276 128538 81540 128548
rect 111996 128604 112260 128614
rect 112052 128548 112100 128604
rect 112156 128548 112204 128604
rect 111996 128538 112260 128548
rect 65916 127820 66180 127830
rect 65972 127764 66020 127820
rect 66076 127764 66124 127820
rect 65916 127754 66180 127764
rect 96636 127820 96900 127830
rect 96692 127764 96740 127820
rect 96796 127764 96844 127820
rect 96636 127754 96900 127764
rect 81276 127036 81540 127046
rect 81332 126980 81380 127036
rect 81436 126980 81484 127036
rect 81276 126970 81540 126980
rect 111996 127036 112260 127046
rect 112052 126980 112100 127036
rect 112156 126980 112204 127036
rect 111996 126970 112260 126980
rect 118076 126754 118132 126766
rect 118076 126702 118078 126754
rect 118130 126702 118132 126754
rect 118076 126420 118132 126702
rect 118076 126354 118132 126364
rect 65916 126252 66180 126262
rect 65972 126196 66020 126252
rect 66076 126196 66124 126252
rect 65916 126186 66180 126196
rect 96636 126252 96900 126262
rect 96692 126196 96740 126252
rect 96796 126196 96844 126252
rect 96636 126186 96900 126196
rect 81276 125468 81540 125478
rect 81332 125412 81380 125468
rect 81436 125412 81484 125468
rect 81276 125402 81540 125412
rect 111996 125468 112260 125478
rect 112052 125412 112100 125468
rect 112156 125412 112204 125468
rect 111996 125402 112260 125412
rect 65916 124684 66180 124694
rect 65972 124628 66020 124684
rect 66076 124628 66124 124684
rect 65916 124618 66180 124628
rect 96636 124684 96900 124694
rect 96692 124628 96740 124684
rect 96796 124628 96844 124684
rect 96636 124618 96900 124628
rect 118076 124066 118132 124078
rect 118076 124014 118078 124066
rect 118130 124014 118132 124066
rect 81276 123900 81540 123910
rect 81332 123844 81380 123900
rect 81436 123844 81484 123900
rect 81276 123834 81540 123844
rect 111996 123900 112260 123910
rect 112052 123844 112100 123900
rect 112156 123844 112204 123900
rect 111996 123834 112260 123844
rect 118076 123732 118132 124014
rect 118076 123666 118132 123676
rect 65916 123116 66180 123126
rect 65972 123060 66020 123116
rect 66076 123060 66124 123116
rect 65916 123050 66180 123060
rect 96636 123116 96900 123126
rect 96692 123060 96740 123116
rect 96796 123060 96844 123116
rect 96636 123050 96900 123060
rect 81276 122332 81540 122342
rect 81332 122276 81380 122332
rect 81436 122276 81484 122332
rect 81276 122266 81540 122276
rect 111996 122332 112260 122342
rect 112052 122276 112100 122332
rect 112156 122276 112204 122332
rect 111996 122266 112260 122276
rect 65916 121548 66180 121558
rect 65972 121492 66020 121548
rect 66076 121492 66124 121548
rect 65916 121482 66180 121492
rect 96636 121548 96900 121558
rect 96692 121492 96740 121548
rect 96796 121492 96844 121548
rect 96636 121482 96900 121492
rect 81276 120764 81540 120774
rect 81332 120708 81380 120764
rect 81436 120708 81484 120764
rect 81276 120698 81540 120708
rect 111996 120764 112260 120774
rect 112052 120708 112100 120764
rect 112156 120708 112204 120764
rect 111996 120698 112260 120708
rect 65916 119980 66180 119990
rect 65972 119924 66020 119980
rect 66076 119924 66124 119980
rect 65916 119914 66180 119924
rect 96636 119980 96900 119990
rect 96692 119924 96740 119980
rect 96796 119924 96844 119980
rect 96636 119914 96900 119924
rect 81276 119196 81540 119206
rect 81332 119140 81380 119196
rect 81436 119140 81484 119196
rect 81276 119130 81540 119140
rect 111996 119196 112260 119206
rect 112052 119140 112100 119196
rect 112156 119140 112204 119196
rect 111996 119130 112260 119140
rect 65916 118412 66180 118422
rect 65972 118356 66020 118412
rect 66076 118356 66124 118412
rect 65916 118346 66180 118356
rect 96636 118412 96900 118422
rect 96692 118356 96740 118412
rect 96796 118356 96844 118412
rect 96636 118346 96900 118356
rect 81276 117628 81540 117638
rect 81332 117572 81380 117628
rect 81436 117572 81484 117628
rect 81276 117562 81540 117572
rect 111996 117628 112260 117638
rect 112052 117572 112100 117628
rect 112156 117572 112204 117628
rect 111996 117562 112260 117572
rect 65916 116844 66180 116854
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 65916 116778 66180 116788
rect 96636 116844 96900 116854
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96636 116778 96900 116788
rect 118076 116340 118132 116350
rect 118076 116246 118132 116284
rect 81276 116060 81540 116070
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81276 115994 81540 116004
rect 111996 116060 112260 116070
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 111996 115994 112260 116004
rect 118076 115778 118132 115790
rect 118076 115726 118078 115778
rect 118130 115726 118132 115778
rect 65916 115276 66180 115286
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 65916 115210 66180 115220
rect 96636 115276 96900 115286
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96636 115210 96900 115220
rect 118076 114996 118132 115726
rect 118076 114930 118132 114940
rect 81276 114492 81540 114502
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81276 114426 81540 114436
rect 111996 114492 112260 114502
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 111996 114426 112260 114436
rect 118076 114324 118132 114334
rect 117628 114322 118132 114324
rect 117628 114270 118078 114322
rect 118130 114270 118132 114322
rect 117628 114268 118132 114270
rect 65916 113708 66180 113718
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 65916 113642 66180 113652
rect 96636 113708 96900 113718
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96636 113642 96900 113652
rect 117628 113652 117684 114268
rect 118076 114258 118132 114268
rect 117628 113586 117684 113596
rect 81276 112924 81540 112934
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81276 112858 81540 112868
rect 111996 112924 112260 112934
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 111996 112858 112260 112868
rect 65916 112140 66180 112150
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 65916 112074 66180 112084
rect 96636 112140 96900 112150
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96636 112074 96900 112084
rect 118076 111636 118132 111646
rect 118076 111542 118132 111580
rect 81276 111356 81540 111366
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81276 111290 81540 111300
rect 111996 111356 112260 111366
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 111996 111290 112260 111300
rect 118076 111074 118132 111086
rect 118076 111022 118078 111074
rect 118130 111022 118132 111074
rect 65916 110572 66180 110582
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 65916 110506 66180 110516
rect 96636 110572 96900 110582
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96636 110506 96900 110516
rect 118076 110292 118132 111022
rect 118076 110226 118132 110236
rect 81276 109788 81540 109798
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81276 109722 81540 109732
rect 111996 109788 112260 109798
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 111996 109722 112260 109732
rect 65916 109004 66180 109014
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 65916 108938 66180 108948
rect 96636 109004 96900 109014
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96636 108938 96900 108948
rect 81276 108220 81540 108230
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81276 108154 81540 108164
rect 111996 108220 112260 108230
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 111996 108154 112260 108164
rect 118076 107938 118132 107950
rect 118076 107886 118078 107938
rect 118130 107886 118132 107938
rect 118076 107604 118132 107886
rect 118076 107538 118132 107548
rect 65916 107436 66180 107446
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 65916 107370 66180 107380
rect 96636 107436 96900 107446
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96636 107370 96900 107380
rect 118076 106818 118132 106830
rect 118076 106766 118078 106818
rect 118130 106766 118132 106818
rect 81276 106652 81540 106662
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81276 106586 81540 106596
rect 111996 106652 112260 106662
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 111996 106586 112260 106596
rect 118076 106260 118132 106766
rect 118076 106194 118132 106204
rect 65916 105868 66180 105878
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 65916 105802 66180 105812
rect 96636 105868 96900 105878
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96636 105802 96900 105812
rect 81276 105084 81540 105094
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81276 105018 81540 105028
rect 111996 105084 112260 105094
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 111996 105018 112260 105028
rect 65916 104300 66180 104310
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 65916 104234 66180 104244
rect 96636 104300 96900 104310
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96636 104234 96900 104244
rect 81276 103516 81540 103526
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81276 103450 81540 103460
rect 111996 103516 112260 103526
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 111996 103450 112260 103460
rect 118076 103234 118132 103246
rect 118076 103182 118078 103234
rect 118130 103182 118132 103234
rect 118076 102900 118132 103182
rect 118076 102834 118132 102844
rect 65916 102732 66180 102742
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 65916 102666 66180 102676
rect 96636 102732 96900 102742
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96636 102666 96900 102676
rect 81276 101948 81540 101958
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81276 101882 81540 101892
rect 111996 101948 112260 101958
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 111996 101882 112260 101892
rect 65916 101164 66180 101174
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 65916 101098 66180 101108
rect 96636 101164 96900 101174
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96636 101098 96900 101108
rect 81276 100380 81540 100390
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81276 100314 81540 100324
rect 111996 100380 112260 100390
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 111996 100314 112260 100324
rect 65916 99596 66180 99606
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 65916 99530 66180 99540
rect 96636 99596 96900 99606
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96636 99530 96900 99540
rect 81276 98812 81540 98822
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81276 98746 81540 98756
rect 111996 98812 112260 98822
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 111996 98746 112260 98756
rect 118076 98530 118132 98542
rect 118076 98478 118078 98530
rect 118130 98478 118132 98530
rect 118076 98196 118132 98478
rect 118076 98130 118132 98140
rect 65916 98028 66180 98038
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 65916 97962 66180 97972
rect 96636 98028 96900 98038
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96636 97962 96900 97972
rect 118076 97410 118132 97422
rect 118076 97358 118078 97410
rect 118130 97358 118132 97410
rect 81276 97244 81540 97254
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81276 97178 81540 97188
rect 111996 97244 112260 97254
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 111996 97178 112260 97188
rect 118076 96852 118132 97358
rect 118076 96786 118132 96796
rect 65916 96460 66180 96470
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 65916 96394 66180 96404
rect 96636 96460 96900 96470
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96636 96394 96900 96404
rect 118076 95842 118132 95854
rect 118076 95790 118078 95842
rect 118130 95790 118132 95842
rect 81276 95676 81540 95686
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81276 95610 81540 95620
rect 111996 95676 112260 95686
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 111996 95610 112260 95620
rect 118076 95508 118132 95790
rect 118076 95442 118132 95452
rect 65916 94892 66180 94902
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 65916 94826 66180 94836
rect 96636 94892 96900 94902
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96636 94826 96900 94836
rect 81276 94108 81540 94118
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81276 94042 81540 94052
rect 111996 94108 112260 94118
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 111996 94042 112260 94052
rect 65916 93324 66180 93334
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 65916 93258 66180 93268
rect 96636 93324 96900 93334
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96636 93258 96900 93268
rect 81276 92540 81540 92550
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81276 92474 81540 92484
rect 111996 92540 112260 92550
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 111996 92474 112260 92484
rect 65916 91756 66180 91766
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 65916 91690 66180 91700
rect 96636 91756 96900 91766
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96636 91690 96900 91700
rect 118076 91138 118132 91150
rect 118076 91086 118078 91138
rect 118130 91086 118132 91138
rect 81276 90972 81540 90982
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81276 90906 81540 90916
rect 111996 90972 112260 90982
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 111996 90906 112260 90916
rect 118076 90804 118132 91086
rect 118076 90738 118132 90748
rect 65916 90188 66180 90198
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 65916 90122 66180 90132
rect 96636 90188 96900 90198
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96636 90122 96900 90132
rect 81276 89404 81540 89414
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81276 89338 81540 89348
rect 111996 89404 112260 89414
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 111996 89338 112260 89348
rect 65916 88620 66180 88630
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 65916 88554 66180 88564
rect 96636 88620 96900 88630
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96636 88554 96900 88564
rect 118076 88116 118132 88126
rect 118076 88022 118132 88060
rect 81276 87836 81540 87846
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81276 87770 81540 87780
rect 111996 87836 112260 87846
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 111996 87770 112260 87780
rect 65916 87052 66180 87062
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 65916 86986 66180 86996
rect 96636 87052 96900 87062
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96636 86986 96900 86996
rect 81276 86268 81540 86278
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81276 86202 81540 86212
rect 111996 86268 112260 86278
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 111996 86202 112260 86212
rect 65916 85484 66180 85494
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 65916 85418 66180 85428
rect 96636 85484 96900 85494
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96636 85418 96900 85428
rect 81276 84700 81540 84710
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81276 84634 81540 84644
rect 111996 84700 112260 84710
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 111996 84634 112260 84644
rect 118076 84418 118132 84430
rect 118076 84366 118078 84418
rect 118130 84366 118132 84418
rect 118076 84084 118132 84366
rect 118076 84018 118132 84028
rect 65916 83916 66180 83926
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 65916 83850 66180 83860
rect 96636 83916 96900 83926
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96636 83850 96900 83860
rect 81276 83132 81540 83142
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81276 83066 81540 83076
rect 111996 83132 112260 83142
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 111996 83066 112260 83076
rect 118076 82850 118132 82862
rect 118076 82798 118078 82850
rect 118130 82798 118132 82850
rect 65916 82348 66180 82358
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 65916 82282 66180 82292
rect 96636 82348 96900 82358
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96636 82282 96900 82292
rect 118076 82068 118132 82798
rect 118076 82002 118132 82012
rect 81276 81564 81540 81574
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81276 81498 81540 81508
rect 111996 81564 112260 81574
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 111996 81498 112260 81508
rect 65916 80780 66180 80790
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 65916 80714 66180 80724
rect 96636 80780 96900 80790
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96636 80714 96900 80724
rect 81276 79996 81540 80006
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81276 79930 81540 79940
rect 111996 79996 112260 80006
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 111996 79930 112260 79940
rect 118076 79714 118132 79726
rect 118076 79662 118078 79714
rect 118130 79662 118132 79714
rect 118076 79380 118132 79662
rect 118076 79314 118132 79324
rect 65916 79212 66180 79222
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 65916 79146 66180 79156
rect 96636 79212 96900 79222
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96636 79146 96900 79156
rect 81276 78428 81540 78438
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81276 78362 81540 78372
rect 111996 78428 112260 78438
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 111996 78362 112260 78372
rect 65916 77644 66180 77654
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 65916 77578 66180 77588
rect 96636 77644 96900 77654
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96636 77578 96900 77588
rect 118076 77026 118132 77038
rect 118076 76974 118078 77026
rect 118130 76974 118132 77026
rect 81276 76860 81540 76870
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81276 76794 81540 76804
rect 111996 76860 112260 76870
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 111996 76794 112260 76804
rect 118076 76692 118132 76974
rect 118076 76626 118132 76636
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 96636 76076 96900 76086
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96636 76010 96900 76020
rect 81276 75292 81540 75302
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81276 75226 81540 75236
rect 111996 75292 112260 75302
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 111996 75226 112260 75236
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 96636 74508 96900 74518
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96636 74442 96900 74452
rect 118076 73890 118132 73902
rect 118076 73838 118078 73890
rect 118130 73838 118132 73890
rect 81276 73724 81540 73734
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81276 73658 81540 73668
rect 111996 73724 112260 73734
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 111996 73658 112260 73668
rect 118076 73332 118132 73838
rect 118076 73266 118132 73276
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 96636 72940 96900 72950
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96636 72874 96900 72884
rect 81276 72156 81540 72166
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81276 72090 81540 72100
rect 111996 72156 112260 72166
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 111996 72090 112260 72100
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 96636 71372 96900 71382
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96636 71306 96900 71316
rect 81276 70588 81540 70598
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81276 70522 81540 70532
rect 111996 70588 112260 70598
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 111996 70522 112260 70532
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 96636 69804 96900 69814
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96636 69738 96900 69748
rect 118076 69300 118132 69310
rect 118076 69206 118132 69244
rect 81276 69020 81540 69030
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81276 68954 81540 68964
rect 111996 69020 112260 69030
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 111996 68954 112260 68964
rect 118076 68738 118132 68750
rect 118076 68686 118078 68738
rect 118130 68686 118132 68738
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 96636 68236 96900 68246
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96636 68170 96900 68180
rect 60620 67890 60676 67900
rect 118076 67956 118132 68686
rect 118076 67890 118132 67900
rect 59612 67790 59614 67842
rect 59666 67790 59668 67842
rect 59612 67778 59668 67790
rect 59276 67618 59332 67630
rect 59276 67566 59278 67618
rect 59330 67566 59332 67618
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 4060 45266 4116 45276
rect 2604 45042 2660 45052
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 2268 40898 2324 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 1820 40338 1876 40348
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 1820 39394 1876 39406
rect 1820 39342 1822 39394
rect 1874 39342 1876 39394
rect 1820 39060 1876 39342
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 1820 38994 1876 39004
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 1820 37378 1876 37390
rect 1820 37326 1822 37378
rect 1874 37326 1876 37378
rect 1820 37044 1876 37326
rect 1820 36978 1876 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1820 36258 1876 36270
rect 1820 36206 1822 36258
rect 1874 36206 1876 36258
rect 1820 35700 1876 36206
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 1820 35634 1876 35644
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 1820 33122 1876 33134
rect 1820 33070 1822 33122
rect 1874 33070 1876 33122
rect 1820 33012 1876 33070
rect 1820 32946 1876 32956
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 1820 29986 1876 29998
rect 1820 29934 1822 29986
rect 1874 29934 1876 29986
rect 1820 29652 1876 29934
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 1820 29586 1876 29596
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 1820 26402 1876 26414
rect 1820 26350 1822 26402
rect 1874 26350 1876 26402
rect 1820 25620 1876 26350
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 1820 25554 1876 25564
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 1820 23266 1876 23278
rect 1820 23214 1822 23266
rect 1874 23214 1876 23266
rect 1820 22932 1876 23214
rect 1820 22866 1876 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 1820 21698 1876 21710
rect 1820 21646 1822 21698
rect 1874 21646 1876 21698
rect 1820 20916 1876 21646
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1820 20850 1876 20860
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 1820 18562 1876 18574
rect 1820 18510 1822 18562
rect 1874 18510 1876 18562
rect 1820 18228 1876 18510
rect 1820 18162 1876 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1820 17442 1876 17454
rect 1820 17390 1822 17442
rect 1874 17390 1876 17442
rect 1820 16884 1876 17390
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 1820 16818 1876 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 1820 11170 1876 11182
rect 1820 11118 1822 11170
rect 1874 11118 1876 11170
rect 1820 10836 1876 11118
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 1820 10770 1876 10780
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 1820 8034 1876 8046
rect 1820 7982 1822 8034
rect 1874 7982 1876 8034
rect 1820 7476 1876 7982
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 1820 7410 1876 7420
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 1820 6466 1876 6478
rect 1820 6414 1822 6466
rect 1874 6414 1876 6466
rect 1820 6132 1876 6414
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 1820 6066 1876 6076
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 1820 4898 1876 4910
rect 1820 4846 1822 4898
rect 1874 4846 1876 4898
rect 1820 4788 1876 4846
rect 1820 4722 1876 4732
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 1820 4450 1876 4462
rect 1820 4398 1822 4450
rect 1874 4398 1876 4450
rect 28 2324 84 2334
rect 28 800 84 2268
rect 1820 2324 1876 4398
rect 20636 4228 20692 66780
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 59276 48132 59332 67566
rect 118076 67618 118132 67630
rect 118076 67566 118078 67618
rect 118130 67566 118132 67618
rect 81276 67452 81540 67462
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81276 67386 81540 67396
rect 111996 67452 112260 67462
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 111996 67386 112260 67396
rect 118076 67284 118132 67566
rect 118076 67218 118132 67228
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 96636 66668 96900 66678
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96636 66602 96900 66612
rect 81276 65884 81540 65894
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81276 65818 81540 65828
rect 111996 65884 112260 65894
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 111996 65818 112260 65828
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 96636 65100 96900 65110
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96636 65034 96900 65044
rect 81276 64316 81540 64326
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81276 64250 81540 64260
rect 111996 64316 112260 64326
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 111996 64250 112260 64260
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 96636 63532 96900 63542
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96636 63466 96900 63476
rect 81276 62748 81540 62758
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81276 62682 81540 62692
rect 111996 62748 112260 62758
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 111996 62682 112260 62692
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 96636 61964 96900 61974
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96636 61898 96900 61908
rect 81276 61180 81540 61190
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81276 61114 81540 61124
rect 111996 61180 112260 61190
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 111996 61114 112260 61124
rect 118076 60898 118132 60910
rect 118076 60846 118078 60898
rect 118130 60846 118132 60898
rect 118076 60564 118132 60846
rect 118076 60498 118132 60508
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 96636 60396 96900 60406
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96636 60330 96900 60340
rect 118076 59892 118132 59902
rect 118076 59798 118132 59836
rect 81276 59612 81540 59622
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81276 59546 81540 59556
rect 111996 59612 112260 59622
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 111996 59546 112260 59556
rect 118076 59330 118132 59342
rect 118076 59278 118078 59330
rect 118130 59278 118132 59330
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 96636 58828 96900 58838
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96636 58762 96900 58772
rect 118076 58548 118132 59278
rect 118076 58482 118132 58492
rect 81276 58044 81540 58054
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81276 57978 81540 57988
rect 111996 58044 112260 58054
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 111996 57978 112260 57988
rect 118076 57762 118132 57774
rect 118076 57710 118078 57762
rect 118130 57710 118132 57762
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 96636 57260 96900 57270
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96636 57194 96900 57204
rect 118076 57204 118132 57710
rect 118076 57138 118132 57148
rect 81276 56476 81540 56486
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81276 56410 81540 56420
rect 111996 56476 112260 56486
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 111996 56410 112260 56420
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 96636 55692 96900 55702
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96636 55626 96900 55636
rect 81276 54908 81540 54918
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81276 54842 81540 54852
rect 111996 54908 112260 54918
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 111996 54842 112260 54852
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 96636 54124 96900 54134
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96636 54058 96900 54068
rect 118076 53506 118132 53518
rect 118076 53454 118078 53506
rect 118130 53454 118132 53506
rect 81276 53340 81540 53350
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81276 53274 81540 53284
rect 111996 53340 112260 53350
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 111996 53274 112260 53284
rect 118076 53284 118132 53454
rect 118076 53218 118132 53228
rect 118076 53058 118132 53070
rect 118076 53006 118078 53058
rect 118130 53006 118132 53058
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 96636 52556 96900 52566
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96636 52490 96900 52500
rect 118076 52500 118132 53006
rect 118076 52434 118132 52444
rect 81276 51772 81540 51782
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81276 51706 81540 51716
rect 111996 51772 112260 51782
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 111996 51706 112260 51716
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 96636 50988 96900 50998
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96636 50922 96900 50932
rect 81276 50204 81540 50214
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81276 50138 81540 50148
rect 111996 50204 112260 50214
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 111996 50138 112260 50148
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 96636 49420 96900 49430
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96636 49354 96900 49364
rect 81276 48636 81540 48646
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81276 48570 81540 48580
rect 111996 48636 112260 48646
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 111996 48570 112260 48580
rect 59276 48066 59332 48076
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 96636 47852 96900 47862
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96636 47786 96900 47796
rect 118076 47234 118132 47246
rect 118076 47182 118078 47234
rect 118130 47182 118132 47234
rect 118076 47124 118132 47182
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 81276 47068 81540 47078
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81276 47002 81540 47012
rect 111996 47068 112260 47078
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 118076 47058 118132 47068
rect 111996 47002 112260 47012
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 96636 46284 96900 46294
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96636 46218 96900 46228
rect 118076 45666 118132 45678
rect 118076 45614 118078 45666
rect 118130 45614 118132 45666
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 81276 45500 81540 45510
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81276 45434 81540 45444
rect 111996 45500 112260 45510
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 111996 45434 112260 45444
rect 118076 45108 118132 45614
rect 118076 45042 118132 45052
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 96636 44716 96900 44726
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96636 44650 96900 44660
rect 118076 44098 118132 44110
rect 118076 44046 118078 44098
rect 118130 44046 118132 44098
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 81276 43932 81540 43942
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81276 43866 81540 43876
rect 111996 43932 112260 43942
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 111996 43866 112260 43876
rect 118076 43764 118132 44046
rect 118076 43698 118132 43708
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 96636 43148 96900 43158
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96636 43082 96900 43092
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 81276 42364 81540 42374
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81276 42298 81540 42308
rect 111996 42364 112260 42374
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 111996 42298 112260 42308
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 96636 41580 96900 41590
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96636 41514 96900 41524
rect 59948 41074 60004 41086
rect 59948 41022 59950 41074
rect 60002 41022 60004 41074
rect 59388 40964 59444 40974
rect 59388 40870 59444 40908
rect 59948 40964 60004 41022
rect 118076 41076 118132 41086
rect 118076 40982 118132 41020
rect 59948 40898 60004 40908
rect 60284 40962 60340 40974
rect 60284 40910 60286 40962
rect 60338 40910 60340 40962
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 60284 35588 60340 40910
rect 81276 40796 81540 40806
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81276 40730 81540 40740
rect 111996 40796 112260 40806
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 111996 40730 112260 40740
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 96636 40012 96900 40022
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96636 39946 96900 39956
rect 81276 39228 81540 39238
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81276 39162 81540 39172
rect 111996 39228 112260 39238
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 111996 39162 112260 39172
rect 118076 38946 118132 38958
rect 118076 38894 118078 38946
rect 118130 38894 118132 38946
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 96636 38444 96900 38454
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96636 38378 96900 38388
rect 118076 38388 118132 38894
rect 118076 38322 118132 38332
rect 81276 37660 81540 37670
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81276 37594 81540 37604
rect 111996 37660 112260 37670
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 111996 37594 112260 37604
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 96636 36876 96900 36886
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96636 36810 96900 36820
rect 117740 36372 117796 36382
rect 81276 36092 81540 36102
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81276 36026 81540 36036
rect 111996 36092 112260 36102
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 111996 36026 112260 36036
rect 117740 35810 117796 36316
rect 117740 35758 117742 35810
rect 117794 35758 117796 35810
rect 117740 35746 117796 35758
rect 116844 35698 116900 35710
rect 116844 35646 116846 35698
rect 116898 35646 116900 35698
rect 60284 35522 60340 35532
rect 116284 35588 116340 35598
rect 116284 35494 116340 35532
rect 116844 35588 116900 35646
rect 116844 35522 116900 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 96636 35308 96900 35318
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96636 35242 96900 35252
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 81276 34524 81540 34534
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81276 34458 81540 34468
rect 111996 34524 112260 34534
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 111996 34458 112260 34468
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 96636 33740 96900 33750
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96636 33674 96900 33684
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 81276 32956 81540 32966
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81276 32890 81540 32900
rect 111996 32956 112260 32966
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 111996 32890 112260 32900
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 96636 32172 96900 32182
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96636 32106 96900 32116
rect 118076 31554 118132 31566
rect 118076 31502 118078 31554
rect 118130 31502 118132 31554
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 81276 31388 81540 31398
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81276 31322 81540 31332
rect 111996 31388 112260 31398
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 111996 31322 112260 31332
rect 118076 30996 118132 31502
rect 118076 30930 118132 30940
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 96636 30604 96900 30614
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96636 30538 96900 30548
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 81276 29820 81540 29830
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81276 29754 81540 29764
rect 111996 29820 112260 29830
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 111996 29754 112260 29764
rect 118076 29538 118132 29550
rect 118076 29486 118078 29538
rect 118130 29486 118132 29538
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 96636 29036 96900 29046
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96636 28970 96900 28980
rect 118076 28980 118132 29486
rect 118076 28914 118132 28924
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 81276 28252 81540 28262
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81276 28186 81540 28196
rect 111996 28252 112260 28262
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 111996 28186 112260 28196
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 96636 27468 96900 27478
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96636 27402 96900 27412
rect 118076 26850 118132 26862
rect 118076 26798 118078 26850
rect 118130 26798 118132 26850
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 81276 26684 81540 26694
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81276 26618 81540 26628
rect 111996 26684 112260 26694
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 111996 26618 112260 26628
rect 118076 26292 118132 26798
rect 118076 26226 118132 26236
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 96636 25900 96900 25910
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96636 25834 96900 25844
rect 118076 25282 118132 25294
rect 118076 25230 118078 25282
rect 118130 25230 118132 25282
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 81276 25116 81540 25126
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81276 25050 81540 25060
rect 111996 25116 112260 25126
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 111996 25050 112260 25060
rect 118076 24948 118132 25230
rect 118076 24882 118132 24892
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 96636 24332 96900 24342
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96636 24266 96900 24276
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 81276 23548 81540 23558
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81276 23482 81540 23492
rect 111996 23548 112260 23558
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 111996 23482 112260 23492
rect 118076 23266 118132 23278
rect 118076 23214 118078 23266
rect 118130 23214 118132 23266
rect 118076 22932 118132 23214
rect 118076 22866 118132 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 96636 22764 96900 22774
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96636 22698 96900 22708
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 81276 21980 81540 21990
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81276 21914 81540 21924
rect 111996 21980 112260 21990
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 111996 21914 112260 21924
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 96636 21196 96900 21206
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96636 21130 96900 21140
rect 118076 20578 118132 20590
rect 118076 20526 118078 20578
rect 118130 20526 118132 20578
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 81276 20412 81540 20422
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81276 20346 81540 20356
rect 111996 20412 112260 20422
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 111996 20346 112260 20356
rect 118076 20244 118132 20526
rect 118076 20178 118132 20188
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 96636 19628 96900 19638
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96636 19562 96900 19572
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 81276 18844 81540 18854
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81276 18778 81540 18788
rect 111996 18844 112260 18854
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 111996 18778 112260 18788
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 96636 18060 96900 18070
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96636 17994 96900 18004
rect 118076 17556 118132 17566
rect 118076 17462 118132 17500
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 81276 17276 81540 17286
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81276 17210 81540 17220
rect 111996 17276 112260 17286
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 111996 17210 112260 17220
rect 118076 16994 118132 17006
rect 118076 16942 118078 16994
rect 118130 16942 118132 16994
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 96636 16492 96900 16502
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96636 16426 96900 16436
rect 118076 16212 118132 16942
rect 118076 16146 118132 16156
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 81276 15708 81540 15718
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81276 15642 81540 15652
rect 111996 15708 112260 15718
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 111996 15642 112260 15652
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 96636 14924 96900 14934
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96636 14858 96900 14868
rect 118076 14306 118132 14318
rect 118076 14254 118078 14306
rect 118130 14254 118132 14306
rect 118076 14196 118132 14254
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 81276 14140 81540 14150
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81276 14074 81540 14084
rect 111996 14140 112260 14150
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 118076 14130 118132 14140
rect 111996 14074 112260 14084
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 96636 13356 96900 13366
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96636 13290 96900 13300
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 81276 12572 81540 12582
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81276 12506 81540 12516
rect 111996 12572 112260 12582
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 111996 12506 112260 12516
rect 118076 12290 118132 12302
rect 118076 12238 118078 12290
rect 118130 12238 118132 12290
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 96636 11788 96900 11798
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96636 11722 96900 11732
rect 118076 11508 118132 12238
rect 118076 11442 118132 11452
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 81276 11004 81540 11014
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81276 10938 81540 10948
rect 111996 11004 112260 11014
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 111996 10938 112260 10948
rect 118076 10722 118132 10734
rect 118076 10670 118078 10722
rect 118130 10670 118132 10722
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 96636 10220 96900 10230
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96636 10154 96900 10164
rect 118076 10164 118132 10670
rect 118076 10098 118132 10108
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 81276 9436 81540 9446
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81276 9370 81540 9380
rect 111996 9436 112260 9446
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 111996 9370 112260 9380
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 96636 8652 96900 8662
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96636 8586 96900 8596
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 81276 7868 81540 7878
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81276 7802 81540 7812
rect 111996 7868 112260 7878
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 111996 7802 112260 7812
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 96636 7084 96900 7094
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96636 7018 96900 7028
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 81276 6300 81540 6310
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81276 6234 81540 6244
rect 111996 6300 112260 6310
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 111996 6234 112260 6244
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 96636 5516 96900 5526
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96636 5450 96900 5460
rect 118076 4900 118132 4910
rect 117964 4898 118132 4900
rect 117964 4846 118078 4898
rect 118130 4846 118132 4898
rect 117964 4844 118132 4846
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 81276 4732 81540 4742
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81276 4666 81540 4676
rect 111996 4732 112260 4742
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 111996 4666 112260 4676
rect 117180 4452 117236 4462
rect 116956 4450 117236 4452
rect 116956 4398 117182 4450
rect 117234 4398 117236 4450
rect 116956 4396 117236 4398
rect 20636 4162 20692 4172
rect 116508 4228 116564 4238
rect 116508 4134 116564 4172
rect 116844 4228 116900 4238
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 96636 3948 96900 3958
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96636 3882 96900 3892
rect 116844 3554 116900 4172
rect 116844 3502 116846 3554
rect 116898 3502 116900 3554
rect 116844 3490 116900 3502
rect 2268 3332 2324 3342
rect 7644 3332 7700 3342
rect 8316 3332 8372 3342
rect 9660 3332 9716 3342
rect 12348 3332 12404 3342
rect 15036 3332 15092 3342
rect 27132 3332 27188 3342
rect 28364 3332 28420 3342
rect 29820 3332 29876 3342
rect 30492 3332 30548 3342
rect 33180 3332 33236 3342
rect 34524 3332 34580 3342
rect 37212 3332 37268 3342
rect 37884 3332 37940 3342
rect 43260 3332 43316 3342
rect 45276 3332 45332 3342
rect 47964 3332 48020 3342
rect 49308 3332 49364 3342
rect 51884 3332 51940 3342
rect 52780 3332 52836 3342
rect 54012 3332 54068 3342
rect 55356 3332 55412 3342
rect 59388 3332 59444 3342
rect 62748 3332 62804 3342
rect 1820 2258 1876 2268
rect 2044 3330 2324 3332
rect 2044 3278 2270 3330
rect 2322 3278 2324 3330
rect 2044 3276 2324 3278
rect 2044 800 2100 3276
rect 2268 3266 2324 3276
rect 7420 3330 7700 3332
rect 7420 3278 7646 3330
rect 7698 3278 7700 3330
rect 7420 3276 7700 3278
rect 7420 800 7476 3276
rect 7644 3266 7700 3276
rect 8092 3330 8372 3332
rect 8092 3278 8318 3330
rect 8370 3278 8372 3330
rect 8092 3276 8372 3278
rect 8092 800 8148 3276
rect 8316 3266 8372 3276
rect 9436 3330 9716 3332
rect 9436 3278 9662 3330
rect 9714 3278 9716 3330
rect 9436 3276 9716 3278
rect 9436 800 9492 3276
rect 9660 3266 9716 3276
rect 12124 3330 12404 3332
rect 12124 3278 12350 3330
rect 12402 3278 12404 3330
rect 12124 3276 12404 3278
rect 12124 800 12180 3276
rect 12348 3266 12404 3276
rect 14812 3330 15092 3332
rect 14812 3278 15038 3330
rect 15090 3278 15092 3330
rect 14812 3276 15092 3278
rect 14812 800 14868 3276
rect 15036 3266 15092 3276
rect 26908 3330 27188 3332
rect 26908 3278 27134 3330
rect 27186 3278 27188 3330
rect 26908 3276 27188 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 26908 800 26964 3276
rect 27132 3266 27188 3276
rect 28252 3330 28420 3332
rect 28252 3278 28366 3330
rect 28418 3278 28420 3330
rect 28252 3276 28420 3278
rect 28252 800 28308 3276
rect 28364 3266 28420 3276
rect 29596 3330 29876 3332
rect 29596 3278 29822 3330
rect 29874 3278 29876 3330
rect 29596 3276 29876 3278
rect 29596 800 29652 3276
rect 29820 3266 29876 3276
rect 30268 3330 30548 3332
rect 30268 3278 30494 3330
rect 30546 3278 30548 3330
rect 30268 3276 30548 3278
rect 30268 800 30324 3276
rect 30492 3266 30548 3276
rect 32956 3330 33236 3332
rect 32956 3278 33182 3330
rect 33234 3278 33236 3330
rect 32956 3276 33236 3278
rect 32956 800 33012 3276
rect 33180 3266 33236 3276
rect 34300 3330 34580 3332
rect 34300 3278 34526 3330
rect 34578 3278 34580 3330
rect 34300 3276 34580 3278
rect 34300 800 34356 3276
rect 34524 3266 34580 3276
rect 36988 3330 37268 3332
rect 36988 3278 37214 3330
rect 37266 3278 37268 3330
rect 36988 3276 37268 3278
rect 36988 800 37044 3276
rect 37212 3266 37268 3276
rect 37660 3330 37940 3332
rect 37660 3278 37886 3330
rect 37938 3278 37940 3330
rect 37660 3276 37940 3278
rect 37660 800 37716 3276
rect 37884 3266 37940 3276
rect 43036 3330 43316 3332
rect 43036 3278 43262 3330
rect 43314 3278 43316 3330
rect 43036 3276 43316 3278
rect 43036 800 43092 3276
rect 43260 3266 43316 3276
rect 45052 3330 45332 3332
rect 45052 3278 45278 3330
rect 45330 3278 45332 3330
rect 45052 3276 45332 3278
rect 45052 800 45108 3276
rect 45276 3266 45332 3276
rect 47740 3330 48020 3332
rect 47740 3278 47966 3330
rect 48018 3278 48020 3330
rect 47740 3276 48020 3278
rect 47740 800 47796 3276
rect 47964 3266 48020 3276
rect 49084 3330 49364 3332
rect 49084 3278 49310 3330
rect 49362 3278 49364 3330
rect 49084 3276 49364 3278
rect 49084 800 49140 3276
rect 49308 3266 49364 3276
rect 51772 3330 51940 3332
rect 51772 3278 51886 3330
rect 51938 3278 51940 3330
rect 51772 3276 51940 3278
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51772 800 51828 3276
rect 51884 3266 51940 3276
rect 52444 3330 52836 3332
rect 52444 3278 52782 3330
rect 52834 3278 52836 3330
rect 52444 3276 52836 3278
rect 52444 800 52500 3276
rect 52780 3266 52836 3276
rect 53788 3330 54068 3332
rect 53788 3278 54014 3330
rect 54066 3278 54068 3330
rect 53788 3276 54068 3278
rect 53788 800 53844 3276
rect 54012 3266 54068 3276
rect 55132 3330 55412 3332
rect 55132 3278 55358 3330
rect 55410 3278 55412 3330
rect 55132 3276 55412 3278
rect 55132 800 55188 3276
rect 55356 3266 55412 3276
rect 59164 3330 59444 3332
rect 59164 3278 59390 3330
rect 59442 3278 59444 3330
rect 59164 3276 59444 3278
rect 59164 800 59220 3276
rect 59388 3266 59444 3276
rect 62524 3330 62804 3332
rect 62524 3278 62750 3330
rect 62802 3278 62804 3330
rect 62524 3276 62804 3278
rect 62524 800 62580 3276
rect 62748 3266 62804 3276
rect 68460 3330 68516 3342
rect 68460 3278 68462 3330
rect 68514 3278 68516 3330
rect 67900 1762 67956 1774
rect 67900 1710 67902 1762
rect 67954 1710 67956 1762
rect 67900 800 67956 1710
rect 68460 1762 68516 3278
rect 68460 1710 68462 1762
rect 68514 1710 68516 1762
rect 68460 1698 68516 1710
rect 68572 3332 68628 3342
rect 68572 800 68628 3276
rect 69132 3332 69188 3342
rect 70140 3332 70196 3342
rect 76300 3332 76356 3342
rect 77532 3332 77588 3342
rect 78876 3332 78932 3342
rect 82908 3332 82964 3342
rect 84924 3332 84980 3342
rect 86268 3332 86324 3342
rect 69132 3238 69188 3276
rect 69916 3330 70196 3332
rect 69916 3278 70142 3330
rect 70194 3278 70196 3330
rect 69916 3276 70196 3278
rect 69916 800 69972 3276
rect 70140 3266 70196 3276
rect 75964 3330 76356 3332
rect 75964 3278 76302 3330
rect 76354 3278 76356 3330
rect 75964 3276 76356 3278
rect 75964 800 76020 3276
rect 76300 3266 76356 3276
rect 77308 3330 77588 3332
rect 77308 3278 77534 3330
rect 77586 3278 77588 3330
rect 77308 3276 77588 3278
rect 77308 800 77364 3276
rect 77532 3266 77588 3276
rect 78652 3330 78932 3332
rect 78652 3278 78878 3330
rect 78930 3278 78932 3330
rect 78652 3276 78932 3278
rect 78652 800 78708 3276
rect 78876 3266 78932 3276
rect 82684 3330 82964 3332
rect 82684 3278 82910 3330
rect 82962 3278 82964 3330
rect 82684 3276 82964 3278
rect 81276 3164 81540 3174
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81276 3098 81540 3108
rect 82684 800 82740 3276
rect 82908 3266 82964 3276
rect 84700 3330 84980 3332
rect 84700 3278 84926 3330
rect 84978 3278 84980 3330
rect 84700 3276 84980 3278
rect 84700 800 84756 3276
rect 84924 3266 84980 3276
rect 86044 3330 86324 3332
rect 86044 3278 86270 3330
rect 86322 3278 86324 3330
rect 86044 3276 86324 3278
rect 86044 800 86100 3276
rect 86268 3266 86324 3276
rect 88060 3330 88116 3342
rect 93660 3332 93716 3342
rect 101052 3332 101108 3342
rect 88060 3278 88062 3330
rect 88114 3278 88116 3330
rect 87388 1874 87444 1886
rect 87388 1822 87390 1874
rect 87442 1822 87444 1874
rect 87388 800 87444 1822
rect 88060 1874 88116 3278
rect 88060 1822 88062 1874
rect 88114 1822 88116 1874
rect 88060 1810 88116 1822
rect 93436 3330 93716 3332
rect 93436 3278 93662 3330
rect 93714 3278 93716 3330
rect 93436 3276 93716 3278
rect 93436 800 93492 3276
rect 93660 3266 93716 3276
rect 100828 3330 101108 3332
rect 100828 3278 101054 3330
rect 101106 3278 101108 3330
rect 100828 3276 101108 3278
rect 100828 800 100884 3276
rect 101052 3266 101108 3276
rect 106876 3332 106932 3342
rect 106876 800 106932 3276
rect 107660 3332 107716 3342
rect 109788 3332 109844 3342
rect 107660 3238 107716 3276
rect 109564 3330 109844 3332
rect 109564 3278 109790 3330
rect 109842 3278 109844 3330
rect 109564 3276 109844 3278
rect 109564 800 109620 3276
rect 109788 3266 109844 3276
rect 111580 3330 111636 3342
rect 111580 3278 111582 3330
rect 111634 3278 111636 3330
rect 110908 1874 110964 1886
rect 110908 1822 110910 1874
rect 110962 1822 110964 1874
rect 110908 800 110964 1822
rect 111580 1874 111636 3278
rect 112476 3330 112532 3342
rect 115836 3332 115892 3342
rect 112476 3278 112478 3330
rect 112530 3278 112532 3330
rect 111996 3164 112260 3174
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 111996 3098 112260 3108
rect 111580 1822 111582 1874
rect 111634 1822 111636 1874
rect 111580 1810 111636 1822
rect 112476 980 112532 3278
rect 112252 924 112532 980
rect 115612 3330 115892 3332
rect 115612 3278 115838 3330
rect 115890 3278 115892 3330
rect 115612 3276 115892 3278
rect 112252 800 112308 924
rect 115612 800 115668 3276
rect 115836 3266 115892 3276
rect 116956 800 117012 4396
rect 117180 4386 117236 4396
rect 117740 3444 117796 3454
rect 117740 3350 117796 3388
rect 0 200 112 800
rect 672 200 784 800
rect 2016 200 2128 800
rect 3360 200 3472 800
rect 4704 200 4816 800
rect 6048 200 6160 800
rect 7392 200 7504 800
rect 8064 200 8176 800
rect 9408 200 9520 800
rect 10752 200 10864 800
rect 12096 200 12208 800
rect 13440 200 13552 800
rect 14784 200 14896 800
rect 15456 200 15568 800
rect 16800 200 16912 800
rect 18144 200 18256 800
rect 19488 200 19600 800
rect 20832 200 20944 800
rect 22176 200 22288 800
rect 22848 200 22960 800
rect 24192 200 24304 800
rect 25536 200 25648 800
rect 26880 200 26992 800
rect 28224 200 28336 800
rect 29568 200 29680 800
rect 30240 200 30352 800
rect 31584 200 31696 800
rect 32928 200 33040 800
rect 34272 200 34384 800
rect 35616 200 35728 800
rect 36960 200 37072 800
rect 37632 200 37744 800
rect 38976 200 39088 800
rect 40320 200 40432 800
rect 41664 200 41776 800
rect 43008 200 43120 800
rect 44352 200 44464 800
rect 45024 200 45136 800
rect 46368 200 46480 800
rect 47712 200 47824 800
rect 49056 200 49168 800
rect 50400 200 50512 800
rect 51744 200 51856 800
rect 52416 200 52528 800
rect 53760 200 53872 800
rect 55104 200 55216 800
rect 56448 200 56560 800
rect 57792 200 57904 800
rect 59136 200 59248 800
rect 59808 200 59920 800
rect 61152 200 61264 800
rect 62496 200 62608 800
rect 63840 200 63952 800
rect 65184 200 65296 800
rect 66528 200 66640 800
rect 67872 200 67984 800
rect 68544 200 68656 800
rect 69888 200 70000 800
rect 71232 200 71344 800
rect 72576 200 72688 800
rect 73920 200 74032 800
rect 75264 200 75376 800
rect 75936 200 76048 800
rect 77280 200 77392 800
rect 78624 200 78736 800
rect 79968 200 80080 800
rect 81312 200 81424 800
rect 82656 200 82768 800
rect 83328 200 83440 800
rect 84672 200 84784 800
rect 86016 200 86128 800
rect 87360 200 87472 800
rect 88704 200 88816 800
rect 90048 200 90160 800
rect 90720 200 90832 800
rect 92064 200 92176 800
rect 93408 200 93520 800
rect 94752 200 94864 800
rect 96096 200 96208 800
rect 97440 200 97552 800
rect 98112 200 98224 800
rect 99456 200 99568 800
rect 100800 200 100912 800
rect 102144 200 102256 800
rect 103488 200 103600 800
rect 104832 200 104944 800
rect 105504 200 105616 800
rect 106848 200 106960 800
rect 108192 200 108304 800
rect 109536 200 109648 800
rect 110880 200 110992 800
rect 112224 200 112336 800
rect 112896 200 113008 800
rect 114240 200 114352 800
rect 115584 200 115696 800
rect 116928 200 117040 800
rect 117964 84 118020 4844
rect 118076 4834 118132 4844
rect 118076 4450 118132 4462
rect 118076 4398 118078 4450
rect 118130 4398 118132 4450
rect 118076 4116 118132 4398
rect 118076 4050 118132 4060
rect 119644 3444 119700 3454
rect 119644 800 119700 3388
rect 118272 200 118384 800
rect 119616 200 119728 800
rect 117964 18 118020 28
<< via2 >>
rect 2492 134428 2548 134484
rect 1820 133084 1876 133140
rect 4476 132522 4532 132524
rect 4476 132470 4478 132522
rect 4478 132470 4530 132522
rect 4530 132470 4532 132522
rect 4476 132468 4532 132470
rect 4580 132522 4636 132524
rect 4580 132470 4582 132522
rect 4582 132470 4634 132522
rect 4634 132470 4636 132522
rect 4580 132468 4636 132470
rect 4684 132522 4740 132524
rect 4684 132470 4686 132522
rect 4686 132470 4738 132522
rect 4738 132470 4740 132522
rect 4684 132468 4740 132470
rect 20188 132188 20244 132244
rect 22092 132242 22148 132244
rect 22092 132190 22094 132242
rect 22094 132190 22146 132242
rect 22146 132190 22148 132242
rect 22092 132188 22148 132190
rect 12796 131964 12852 132020
rect 13580 132018 13636 132020
rect 13580 131966 13582 132018
rect 13582 131966 13634 132018
rect 13634 131966 13636 132018
rect 13580 131964 13636 131966
rect 35196 132522 35252 132524
rect 35196 132470 35198 132522
rect 35198 132470 35250 132522
rect 35250 132470 35252 132522
rect 35196 132468 35252 132470
rect 35300 132522 35356 132524
rect 35300 132470 35302 132522
rect 35302 132470 35354 132522
rect 35354 132470 35356 132522
rect 35300 132468 35356 132470
rect 35404 132522 35460 132524
rect 35404 132470 35406 132522
rect 35406 132470 35458 132522
rect 35458 132470 35460 132522
rect 35404 132468 35460 132470
rect 59836 132076 59892 132132
rect 60844 132130 60900 132132
rect 60844 132078 60846 132130
rect 60846 132078 60898 132130
rect 60898 132078 60900 132130
rect 60844 132076 60900 132078
rect 65916 132522 65972 132524
rect 65916 132470 65918 132522
rect 65918 132470 65970 132522
rect 65970 132470 65972 132522
rect 65916 132468 65972 132470
rect 66020 132522 66076 132524
rect 66020 132470 66022 132522
rect 66022 132470 66074 132522
rect 66074 132470 66076 132522
rect 66020 132468 66076 132470
rect 66124 132522 66180 132524
rect 66124 132470 66126 132522
rect 66126 132470 66178 132522
rect 66178 132470 66180 132522
rect 66124 132468 66180 132470
rect 71932 131964 71988 132020
rect 72380 132018 72436 132020
rect 72380 131966 72382 132018
rect 72382 131966 72434 132018
rect 72434 131966 72436 132018
rect 72380 131964 72436 131966
rect 75292 131964 75348 132020
rect 76300 132018 76356 132020
rect 76300 131966 76302 132018
rect 76302 131966 76354 132018
rect 76354 131966 76356 132018
rect 76300 131964 76356 131966
rect 96636 132522 96692 132524
rect 96636 132470 96638 132522
rect 96638 132470 96690 132522
rect 96690 132470 96692 132522
rect 96636 132468 96692 132470
rect 96740 132522 96796 132524
rect 96740 132470 96742 132522
rect 96742 132470 96794 132522
rect 96794 132470 96796 132522
rect 96740 132468 96796 132470
rect 96844 132522 96900 132524
rect 96844 132470 96846 132522
rect 96846 132470 96898 132522
rect 96898 132470 96900 132522
rect 96844 132468 96900 132470
rect 95452 131964 95508 132020
rect 95900 132018 95956 132020
rect 95900 131966 95902 132018
rect 95902 131966 95954 132018
rect 95954 131966 95956 132018
rect 95900 131964 95956 131966
rect 117292 132412 117348 132468
rect 19836 131738 19892 131740
rect 19836 131686 19838 131738
rect 19838 131686 19890 131738
rect 19890 131686 19892 131738
rect 19836 131684 19892 131686
rect 19940 131738 19996 131740
rect 19940 131686 19942 131738
rect 19942 131686 19994 131738
rect 19994 131686 19996 131738
rect 19940 131684 19996 131686
rect 20044 131738 20100 131740
rect 20044 131686 20046 131738
rect 20046 131686 20098 131738
rect 20098 131686 20100 131738
rect 20044 131684 20100 131686
rect 4476 130954 4532 130956
rect 4476 130902 4478 130954
rect 4478 130902 4530 130954
rect 4530 130902 4532 130954
rect 4476 130900 4532 130902
rect 4580 130954 4636 130956
rect 4580 130902 4582 130954
rect 4582 130902 4634 130954
rect 4634 130902 4636 130954
rect 4580 130900 4636 130902
rect 4684 130954 4740 130956
rect 4684 130902 4686 130954
rect 4686 130902 4738 130954
rect 4738 130902 4740 130954
rect 4684 130900 4740 130902
rect 1820 130450 1876 130452
rect 1820 130398 1822 130450
rect 1822 130398 1874 130450
rect 1874 130398 1876 130450
rect 1820 130396 1876 130398
rect 19836 130170 19892 130172
rect 19836 130118 19838 130170
rect 19838 130118 19890 130170
rect 19890 130118 19892 130170
rect 19836 130116 19892 130118
rect 19940 130170 19996 130172
rect 19940 130118 19942 130170
rect 19942 130118 19994 130170
rect 19994 130118 19996 130170
rect 19940 130116 19996 130118
rect 20044 130170 20100 130172
rect 20044 130118 20046 130170
rect 20046 130118 20098 130170
rect 20098 130118 20100 130170
rect 20044 130116 20100 130118
rect 4476 129386 4532 129388
rect 4476 129334 4478 129386
rect 4478 129334 4530 129386
rect 4530 129334 4532 129386
rect 4476 129332 4532 129334
rect 4580 129386 4636 129388
rect 4580 129334 4582 129386
rect 4582 129334 4634 129386
rect 4634 129334 4636 129386
rect 4580 129332 4636 129334
rect 4684 129386 4740 129388
rect 4684 129334 4686 129386
rect 4686 129334 4738 129386
rect 4738 129334 4740 129386
rect 4684 129332 4740 129334
rect 19836 128602 19892 128604
rect 19836 128550 19838 128602
rect 19838 128550 19890 128602
rect 19890 128550 19892 128602
rect 19836 128548 19892 128550
rect 19940 128602 19996 128604
rect 19940 128550 19942 128602
rect 19942 128550 19994 128602
rect 19994 128550 19996 128602
rect 19940 128548 19996 128550
rect 20044 128602 20100 128604
rect 20044 128550 20046 128602
rect 20046 128550 20098 128602
rect 20098 128550 20100 128602
rect 20044 128548 20100 128550
rect 1820 127708 1876 127764
rect 4476 127818 4532 127820
rect 4476 127766 4478 127818
rect 4478 127766 4530 127818
rect 4530 127766 4532 127818
rect 4476 127764 4532 127766
rect 4580 127818 4636 127820
rect 4580 127766 4582 127818
rect 4582 127766 4634 127818
rect 4634 127766 4636 127818
rect 4580 127764 4636 127766
rect 4684 127818 4740 127820
rect 4684 127766 4686 127818
rect 4686 127766 4738 127818
rect 4738 127766 4740 127818
rect 4684 127764 4740 127766
rect 1820 127036 1876 127092
rect 19836 127034 19892 127036
rect 19836 126982 19838 127034
rect 19838 126982 19890 127034
rect 19890 126982 19892 127034
rect 19836 126980 19892 126982
rect 19940 127034 19996 127036
rect 19940 126982 19942 127034
rect 19942 126982 19994 127034
rect 19994 126982 19996 127034
rect 19940 126980 19996 126982
rect 20044 127034 20100 127036
rect 20044 126982 20046 127034
rect 20046 126982 20098 127034
rect 20098 126982 20100 127034
rect 20044 126980 20100 126982
rect 4476 126250 4532 126252
rect 4476 126198 4478 126250
rect 4478 126198 4530 126250
rect 4530 126198 4532 126250
rect 4476 126196 4532 126198
rect 4580 126250 4636 126252
rect 4580 126198 4582 126250
rect 4582 126198 4634 126250
rect 4634 126198 4636 126250
rect 4580 126196 4636 126198
rect 4684 126250 4740 126252
rect 4684 126198 4686 126250
rect 4686 126198 4738 126250
rect 4738 126198 4740 126250
rect 4684 126196 4740 126198
rect 19836 125466 19892 125468
rect 19836 125414 19838 125466
rect 19838 125414 19890 125466
rect 19890 125414 19892 125466
rect 19836 125412 19892 125414
rect 19940 125466 19996 125468
rect 19940 125414 19942 125466
rect 19942 125414 19994 125466
rect 19994 125414 19996 125466
rect 19940 125412 19996 125414
rect 20044 125466 20100 125468
rect 20044 125414 20046 125466
rect 20046 125414 20098 125466
rect 20098 125414 20100 125466
rect 20044 125412 20100 125414
rect 4476 124682 4532 124684
rect 4476 124630 4478 124682
rect 4478 124630 4530 124682
rect 4530 124630 4532 124682
rect 4476 124628 4532 124630
rect 4580 124682 4636 124684
rect 4580 124630 4582 124682
rect 4582 124630 4634 124682
rect 4634 124630 4636 124682
rect 4580 124628 4636 124630
rect 4684 124682 4740 124684
rect 4684 124630 4686 124682
rect 4686 124630 4738 124682
rect 4738 124630 4740 124682
rect 4684 124628 4740 124630
rect 1820 124348 1876 124404
rect 19836 123898 19892 123900
rect 19836 123846 19838 123898
rect 19838 123846 19890 123898
rect 19890 123846 19892 123898
rect 19836 123844 19892 123846
rect 19940 123898 19996 123900
rect 19940 123846 19942 123898
rect 19942 123846 19994 123898
rect 19994 123846 19996 123898
rect 19940 123844 19996 123846
rect 20044 123898 20100 123900
rect 20044 123846 20046 123898
rect 20046 123846 20098 123898
rect 20098 123846 20100 123898
rect 20044 123844 20100 123846
rect 1820 123004 1876 123060
rect 4476 123114 4532 123116
rect 4476 123062 4478 123114
rect 4478 123062 4530 123114
rect 4530 123062 4532 123114
rect 4476 123060 4532 123062
rect 4580 123114 4636 123116
rect 4580 123062 4582 123114
rect 4582 123062 4634 123114
rect 4634 123062 4636 123114
rect 4580 123060 4636 123062
rect 4684 123114 4740 123116
rect 4684 123062 4686 123114
rect 4686 123062 4738 123114
rect 4738 123062 4740 123114
rect 4684 123060 4740 123062
rect 19836 122330 19892 122332
rect 19836 122278 19838 122330
rect 19838 122278 19890 122330
rect 19890 122278 19892 122330
rect 19836 122276 19892 122278
rect 19940 122330 19996 122332
rect 19940 122278 19942 122330
rect 19942 122278 19994 122330
rect 19994 122278 19996 122330
rect 19940 122276 19996 122278
rect 20044 122330 20100 122332
rect 20044 122278 20046 122330
rect 20046 122278 20098 122330
rect 20098 122278 20100 122330
rect 20044 122276 20100 122278
rect 1820 121660 1876 121716
rect 4476 121546 4532 121548
rect 4476 121494 4478 121546
rect 4478 121494 4530 121546
rect 4530 121494 4532 121546
rect 4476 121492 4532 121494
rect 4580 121546 4636 121548
rect 4580 121494 4582 121546
rect 4582 121494 4634 121546
rect 4634 121494 4636 121546
rect 4580 121492 4636 121494
rect 4684 121546 4740 121548
rect 4684 121494 4686 121546
rect 4686 121494 4738 121546
rect 4738 121494 4740 121546
rect 4684 121492 4740 121494
rect 19836 120762 19892 120764
rect 19836 120710 19838 120762
rect 19838 120710 19890 120762
rect 19890 120710 19892 120762
rect 19836 120708 19892 120710
rect 19940 120762 19996 120764
rect 19940 120710 19942 120762
rect 19942 120710 19994 120762
rect 19994 120710 19996 120762
rect 19940 120708 19996 120710
rect 20044 120762 20100 120764
rect 20044 120710 20046 120762
rect 20046 120710 20098 120762
rect 20098 120710 20100 120762
rect 20044 120708 20100 120710
rect 4476 119978 4532 119980
rect 4476 119926 4478 119978
rect 4478 119926 4530 119978
rect 4530 119926 4532 119978
rect 4476 119924 4532 119926
rect 4580 119978 4636 119980
rect 4580 119926 4582 119978
rect 4582 119926 4634 119978
rect 4634 119926 4636 119978
rect 4580 119924 4636 119926
rect 4684 119978 4740 119980
rect 4684 119926 4686 119978
rect 4686 119926 4738 119978
rect 4738 119926 4740 119978
rect 4684 119924 4740 119926
rect 19836 119194 19892 119196
rect 19836 119142 19838 119194
rect 19838 119142 19890 119194
rect 19890 119142 19892 119194
rect 19836 119140 19892 119142
rect 19940 119194 19996 119196
rect 19940 119142 19942 119194
rect 19942 119142 19994 119194
rect 19994 119142 19996 119194
rect 19940 119140 19996 119142
rect 20044 119194 20100 119196
rect 20044 119142 20046 119194
rect 20046 119142 20098 119194
rect 20098 119142 20100 119194
rect 20044 119140 20100 119142
rect 4476 118410 4532 118412
rect 4476 118358 4478 118410
rect 4478 118358 4530 118410
rect 4530 118358 4532 118410
rect 4476 118356 4532 118358
rect 4580 118410 4636 118412
rect 4580 118358 4582 118410
rect 4582 118358 4634 118410
rect 4634 118358 4636 118410
rect 4580 118356 4636 118358
rect 4684 118410 4740 118412
rect 4684 118358 4686 118410
rect 4686 118358 4738 118410
rect 4738 118358 4740 118410
rect 4684 118356 4740 118358
rect 19836 117626 19892 117628
rect 19836 117574 19838 117626
rect 19838 117574 19890 117626
rect 19890 117574 19892 117626
rect 19836 117572 19892 117574
rect 19940 117626 19996 117628
rect 19940 117574 19942 117626
rect 19942 117574 19994 117626
rect 19994 117574 19996 117626
rect 19940 117572 19996 117574
rect 20044 117626 20100 117628
rect 20044 117574 20046 117626
rect 20046 117574 20098 117626
rect 20098 117574 20100 117626
rect 20044 117572 20100 117574
rect 1820 116956 1876 117012
rect 4476 116842 4532 116844
rect 4476 116790 4478 116842
rect 4478 116790 4530 116842
rect 4530 116790 4532 116842
rect 4476 116788 4532 116790
rect 4580 116842 4636 116844
rect 4580 116790 4582 116842
rect 4582 116790 4634 116842
rect 4634 116790 4636 116842
rect 4580 116788 4636 116790
rect 4684 116842 4740 116844
rect 4684 116790 4686 116842
rect 4686 116790 4738 116842
rect 4738 116790 4740 116842
rect 4684 116788 4740 116790
rect 19836 116058 19892 116060
rect 19836 116006 19838 116058
rect 19838 116006 19890 116058
rect 19890 116006 19892 116058
rect 19836 116004 19892 116006
rect 19940 116058 19996 116060
rect 19940 116006 19942 116058
rect 19942 116006 19994 116058
rect 19994 116006 19996 116058
rect 19940 116004 19996 116006
rect 20044 116058 20100 116060
rect 20044 116006 20046 116058
rect 20046 116006 20098 116058
rect 20098 116006 20100 116058
rect 20044 116004 20100 116006
rect 4476 115274 4532 115276
rect 4476 115222 4478 115274
rect 4478 115222 4530 115274
rect 4530 115222 4532 115274
rect 4476 115220 4532 115222
rect 4580 115274 4636 115276
rect 4580 115222 4582 115274
rect 4582 115222 4634 115274
rect 4634 115222 4636 115274
rect 4580 115220 4636 115222
rect 4684 115274 4740 115276
rect 4684 115222 4686 115274
rect 4686 115222 4738 115274
rect 4738 115222 4740 115274
rect 4684 115220 4740 115222
rect 19836 114490 19892 114492
rect 19836 114438 19838 114490
rect 19838 114438 19890 114490
rect 19890 114438 19892 114490
rect 19836 114436 19892 114438
rect 19940 114490 19996 114492
rect 19940 114438 19942 114490
rect 19942 114438 19994 114490
rect 19994 114438 19996 114490
rect 19940 114436 19996 114438
rect 20044 114490 20100 114492
rect 20044 114438 20046 114490
rect 20046 114438 20098 114490
rect 20098 114438 20100 114490
rect 20044 114436 20100 114438
rect 4476 113706 4532 113708
rect 4476 113654 4478 113706
rect 4478 113654 4530 113706
rect 4530 113654 4532 113706
rect 4476 113652 4532 113654
rect 4580 113706 4636 113708
rect 4580 113654 4582 113706
rect 4582 113654 4634 113706
rect 4634 113654 4636 113706
rect 4580 113652 4636 113654
rect 4684 113706 4740 113708
rect 4684 113654 4686 113706
rect 4686 113654 4738 113706
rect 4738 113654 4740 113706
rect 4684 113652 4740 113654
rect 19836 112922 19892 112924
rect 19836 112870 19838 112922
rect 19838 112870 19890 112922
rect 19890 112870 19892 112922
rect 19836 112868 19892 112870
rect 19940 112922 19996 112924
rect 19940 112870 19942 112922
rect 19942 112870 19994 112922
rect 19994 112870 19996 112922
rect 19940 112868 19996 112870
rect 20044 112922 20100 112924
rect 20044 112870 20046 112922
rect 20046 112870 20098 112922
rect 20098 112870 20100 112922
rect 20044 112868 20100 112870
rect 4476 112138 4532 112140
rect 4476 112086 4478 112138
rect 4478 112086 4530 112138
rect 4530 112086 4532 112138
rect 4476 112084 4532 112086
rect 4580 112138 4636 112140
rect 4580 112086 4582 112138
rect 4582 112086 4634 112138
rect 4634 112086 4636 112138
rect 4580 112084 4636 112086
rect 4684 112138 4740 112140
rect 4684 112086 4686 112138
rect 4686 112086 4738 112138
rect 4738 112086 4740 112138
rect 4684 112084 4740 112086
rect 19836 111354 19892 111356
rect 19836 111302 19838 111354
rect 19838 111302 19890 111354
rect 19890 111302 19892 111354
rect 19836 111300 19892 111302
rect 19940 111354 19996 111356
rect 19940 111302 19942 111354
rect 19942 111302 19994 111354
rect 19994 111302 19996 111354
rect 19940 111300 19996 111302
rect 20044 111354 20100 111356
rect 20044 111302 20046 111354
rect 20046 111302 20098 111354
rect 20098 111302 20100 111354
rect 20044 111300 20100 111302
rect 1820 110908 1876 110964
rect 4476 110570 4532 110572
rect 4476 110518 4478 110570
rect 4478 110518 4530 110570
rect 4530 110518 4532 110570
rect 4476 110516 4532 110518
rect 4580 110570 4636 110572
rect 4580 110518 4582 110570
rect 4582 110518 4634 110570
rect 4634 110518 4636 110570
rect 4580 110516 4636 110518
rect 4684 110570 4740 110572
rect 4684 110518 4686 110570
rect 4686 110518 4738 110570
rect 4738 110518 4740 110570
rect 4684 110516 4740 110518
rect 19836 109786 19892 109788
rect 19836 109734 19838 109786
rect 19838 109734 19890 109786
rect 19890 109734 19892 109786
rect 19836 109732 19892 109734
rect 19940 109786 19996 109788
rect 19940 109734 19942 109786
rect 19942 109734 19994 109786
rect 19994 109734 19996 109786
rect 19940 109732 19996 109734
rect 20044 109786 20100 109788
rect 20044 109734 20046 109786
rect 20046 109734 20098 109786
rect 20098 109734 20100 109786
rect 20044 109732 20100 109734
rect 1820 109564 1876 109620
rect 4476 109002 4532 109004
rect 4476 108950 4478 109002
rect 4478 108950 4530 109002
rect 4530 108950 4532 109002
rect 4476 108948 4532 108950
rect 4580 109002 4636 109004
rect 4580 108950 4582 109002
rect 4582 108950 4634 109002
rect 4634 108950 4636 109002
rect 4580 108948 4636 108950
rect 4684 109002 4740 109004
rect 4684 108950 4686 109002
rect 4686 108950 4738 109002
rect 4738 108950 4740 109002
rect 4684 108948 4740 108950
rect 19836 108218 19892 108220
rect 19836 108166 19838 108218
rect 19838 108166 19890 108218
rect 19890 108166 19892 108218
rect 19836 108164 19892 108166
rect 19940 108218 19996 108220
rect 19940 108166 19942 108218
rect 19942 108166 19994 108218
rect 19994 108166 19996 108218
rect 19940 108164 19996 108166
rect 20044 108218 20100 108220
rect 20044 108166 20046 108218
rect 20046 108166 20098 108218
rect 20098 108166 20100 108218
rect 20044 108164 20100 108166
rect 4476 107434 4532 107436
rect 4476 107382 4478 107434
rect 4478 107382 4530 107434
rect 4530 107382 4532 107434
rect 4476 107380 4532 107382
rect 4580 107434 4636 107436
rect 4580 107382 4582 107434
rect 4582 107382 4634 107434
rect 4634 107382 4636 107434
rect 4580 107380 4636 107382
rect 4684 107434 4740 107436
rect 4684 107382 4686 107434
rect 4686 107382 4738 107434
rect 4738 107382 4740 107434
rect 4684 107380 4740 107382
rect 19836 106650 19892 106652
rect 19836 106598 19838 106650
rect 19838 106598 19890 106650
rect 19890 106598 19892 106650
rect 19836 106596 19892 106598
rect 19940 106650 19996 106652
rect 19940 106598 19942 106650
rect 19942 106598 19994 106650
rect 19994 106598 19996 106650
rect 19940 106596 19996 106598
rect 20044 106650 20100 106652
rect 20044 106598 20046 106650
rect 20046 106598 20098 106650
rect 20098 106598 20100 106650
rect 20044 106596 20100 106598
rect 4476 105866 4532 105868
rect 4476 105814 4478 105866
rect 4478 105814 4530 105866
rect 4530 105814 4532 105866
rect 4476 105812 4532 105814
rect 4580 105866 4636 105868
rect 4580 105814 4582 105866
rect 4582 105814 4634 105866
rect 4634 105814 4636 105866
rect 4580 105812 4636 105814
rect 4684 105866 4740 105868
rect 4684 105814 4686 105866
rect 4686 105814 4738 105866
rect 4738 105814 4740 105866
rect 4684 105812 4740 105814
rect 19836 105082 19892 105084
rect 19836 105030 19838 105082
rect 19838 105030 19890 105082
rect 19890 105030 19892 105082
rect 19836 105028 19892 105030
rect 19940 105082 19996 105084
rect 19940 105030 19942 105082
rect 19942 105030 19994 105082
rect 19994 105030 19996 105082
rect 19940 105028 19996 105030
rect 20044 105082 20100 105084
rect 20044 105030 20046 105082
rect 20046 105030 20098 105082
rect 20098 105030 20100 105082
rect 20044 105028 20100 105030
rect 1820 104860 1876 104916
rect 4476 104298 4532 104300
rect 4476 104246 4478 104298
rect 4478 104246 4530 104298
rect 4530 104246 4532 104298
rect 4476 104244 4532 104246
rect 4580 104298 4636 104300
rect 4580 104246 4582 104298
rect 4582 104246 4634 104298
rect 4634 104246 4636 104298
rect 4580 104244 4636 104246
rect 4684 104298 4740 104300
rect 4684 104246 4686 104298
rect 4686 104246 4738 104298
rect 4738 104246 4740 104298
rect 4684 104244 4740 104246
rect 19836 103514 19892 103516
rect 19836 103462 19838 103514
rect 19838 103462 19890 103514
rect 19890 103462 19892 103514
rect 19836 103460 19892 103462
rect 19940 103514 19996 103516
rect 19940 103462 19942 103514
rect 19942 103462 19994 103514
rect 19994 103462 19996 103514
rect 19940 103460 19996 103462
rect 20044 103514 20100 103516
rect 20044 103462 20046 103514
rect 20046 103462 20098 103514
rect 20098 103462 20100 103514
rect 20044 103460 20100 103462
rect 4476 102730 4532 102732
rect 4476 102678 4478 102730
rect 4478 102678 4530 102730
rect 4530 102678 4532 102730
rect 4476 102676 4532 102678
rect 4580 102730 4636 102732
rect 4580 102678 4582 102730
rect 4582 102678 4634 102730
rect 4634 102678 4636 102730
rect 4580 102676 4636 102678
rect 4684 102730 4740 102732
rect 4684 102678 4686 102730
rect 4686 102678 4738 102730
rect 4738 102678 4740 102730
rect 4684 102676 4740 102678
rect 19836 101946 19892 101948
rect 19836 101894 19838 101946
rect 19838 101894 19890 101946
rect 19890 101894 19892 101946
rect 19836 101892 19892 101894
rect 19940 101946 19996 101948
rect 19940 101894 19942 101946
rect 19942 101894 19994 101946
rect 19994 101894 19996 101946
rect 19940 101892 19996 101894
rect 20044 101946 20100 101948
rect 20044 101894 20046 101946
rect 20046 101894 20098 101946
rect 20098 101894 20100 101946
rect 20044 101892 20100 101894
rect 4476 101162 4532 101164
rect 4476 101110 4478 101162
rect 4478 101110 4530 101162
rect 4530 101110 4532 101162
rect 4476 101108 4532 101110
rect 4580 101162 4636 101164
rect 4580 101110 4582 101162
rect 4582 101110 4634 101162
rect 4634 101110 4636 101162
rect 4580 101108 4636 101110
rect 4684 101162 4740 101164
rect 4684 101110 4686 101162
rect 4686 101110 4738 101162
rect 4738 101110 4740 101162
rect 4684 101108 4740 101110
rect 1820 100828 1876 100884
rect 19836 100378 19892 100380
rect 19836 100326 19838 100378
rect 19838 100326 19890 100378
rect 19890 100326 19892 100378
rect 19836 100324 19892 100326
rect 19940 100378 19996 100380
rect 19940 100326 19942 100378
rect 19942 100326 19994 100378
rect 19994 100326 19996 100378
rect 19940 100324 19996 100326
rect 20044 100378 20100 100380
rect 20044 100326 20046 100378
rect 20046 100326 20098 100378
rect 20098 100326 20100 100378
rect 20044 100324 20100 100326
rect 4476 99594 4532 99596
rect 4476 99542 4478 99594
rect 4478 99542 4530 99594
rect 4530 99542 4532 99594
rect 4476 99540 4532 99542
rect 4580 99594 4636 99596
rect 4580 99542 4582 99594
rect 4582 99542 4634 99594
rect 4634 99542 4636 99594
rect 4580 99540 4636 99542
rect 4684 99594 4740 99596
rect 4684 99542 4686 99594
rect 4686 99542 4738 99594
rect 4738 99542 4740 99594
rect 4684 99540 4740 99542
rect 19836 98810 19892 98812
rect 19836 98758 19838 98810
rect 19838 98758 19890 98810
rect 19890 98758 19892 98810
rect 19836 98756 19892 98758
rect 19940 98810 19996 98812
rect 19940 98758 19942 98810
rect 19942 98758 19994 98810
rect 19994 98758 19996 98810
rect 19940 98756 19996 98758
rect 20044 98810 20100 98812
rect 20044 98758 20046 98810
rect 20046 98758 20098 98810
rect 20098 98758 20100 98810
rect 20044 98756 20100 98758
rect 4476 98026 4532 98028
rect 4476 97974 4478 98026
rect 4478 97974 4530 98026
rect 4530 97974 4532 98026
rect 4476 97972 4532 97974
rect 4580 98026 4636 98028
rect 4580 97974 4582 98026
rect 4582 97974 4634 98026
rect 4634 97974 4636 98026
rect 4580 97972 4636 97974
rect 4684 98026 4740 98028
rect 4684 97974 4686 98026
rect 4686 97974 4738 98026
rect 4738 97974 4740 98026
rect 4684 97972 4740 97974
rect 19836 97242 19892 97244
rect 19836 97190 19838 97242
rect 19838 97190 19890 97242
rect 19890 97190 19892 97242
rect 19836 97188 19892 97190
rect 19940 97242 19996 97244
rect 19940 97190 19942 97242
rect 19942 97190 19994 97242
rect 19994 97190 19996 97242
rect 19940 97188 19996 97190
rect 20044 97242 20100 97244
rect 20044 97190 20046 97242
rect 20046 97190 20098 97242
rect 20098 97190 20100 97242
rect 20044 97188 20100 97190
rect 4476 96458 4532 96460
rect 4476 96406 4478 96458
rect 4478 96406 4530 96458
rect 4530 96406 4532 96458
rect 4476 96404 4532 96406
rect 4580 96458 4636 96460
rect 4580 96406 4582 96458
rect 4582 96406 4634 96458
rect 4634 96406 4636 96458
rect 4580 96404 4636 96406
rect 4684 96458 4740 96460
rect 4684 96406 4686 96458
rect 4686 96406 4738 96458
rect 4738 96406 4740 96458
rect 4684 96404 4740 96406
rect 1820 96124 1876 96180
rect 19836 95674 19892 95676
rect 19836 95622 19838 95674
rect 19838 95622 19890 95674
rect 19890 95622 19892 95674
rect 19836 95620 19892 95622
rect 19940 95674 19996 95676
rect 19940 95622 19942 95674
rect 19942 95622 19994 95674
rect 19994 95622 19996 95674
rect 19940 95620 19996 95622
rect 20044 95674 20100 95676
rect 20044 95622 20046 95674
rect 20046 95622 20098 95674
rect 20098 95622 20100 95674
rect 20044 95620 20100 95622
rect 1820 94780 1876 94836
rect 4476 94890 4532 94892
rect 4476 94838 4478 94890
rect 4478 94838 4530 94890
rect 4530 94838 4532 94890
rect 4476 94836 4532 94838
rect 4580 94890 4636 94892
rect 4580 94838 4582 94890
rect 4582 94838 4634 94890
rect 4634 94838 4636 94890
rect 4580 94836 4636 94838
rect 4684 94890 4740 94892
rect 4684 94838 4686 94890
rect 4686 94838 4738 94890
rect 4738 94838 4740 94890
rect 4684 94836 4740 94838
rect 19836 94106 19892 94108
rect 19836 94054 19838 94106
rect 19838 94054 19890 94106
rect 19890 94054 19892 94106
rect 19836 94052 19892 94054
rect 19940 94106 19996 94108
rect 19940 94054 19942 94106
rect 19942 94054 19994 94106
rect 19994 94054 19996 94106
rect 19940 94052 19996 94054
rect 20044 94106 20100 94108
rect 20044 94054 20046 94106
rect 20046 94054 20098 94106
rect 20098 94054 20100 94106
rect 20044 94052 20100 94054
rect 4476 93322 4532 93324
rect 4476 93270 4478 93322
rect 4478 93270 4530 93322
rect 4530 93270 4532 93322
rect 4476 93268 4532 93270
rect 4580 93322 4636 93324
rect 4580 93270 4582 93322
rect 4582 93270 4634 93322
rect 4634 93270 4636 93322
rect 4580 93268 4636 93270
rect 4684 93322 4740 93324
rect 4684 93270 4686 93322
rect 4686 93270 4738 93322
rect 4738 93270 4740 93322
rect 4684 93268 4740 93270
rect 19836 92538 19892 92540
rect 19836 92486 19838 92538
rect 19838 92486 19890 92538
rect 19890 92486 19892 92538
rect 19836 92484 19892 92486
rect 19940 92538 19996 92540
rect 19940 92486 19942 92538
rect 19942 92486 19994 92538
rect 19994 92486 19996 92538
rect 19940 92484 19996 92486
rect 20044 92538 20100 92540
rect 20044 92486 20046 92538
rect 20046 92486 20098 92538
rect 20098 92486 20100 92538
rect 20044 92484 20100 92486
rect 1820 92092 1876 92148
rect 4476 91754 4532 91756
rect 4476 91702 4478 91754
rect 4478 91702 4530 91754
rect 4530 91702 4532 91754
rect 4476 91700 4532 91702
rect 4580 91754 4636 91756
rect 4580 91702 4582 91754
rect 4582 91702 4634 91754
rect 4634 91702 4636 91754
rect 4580 91700 4636 91702
rect 4684 91754 4740 91756
rect 4684 91702 4686 91754
rect 4686 91702 4738 91754
rect 4738 91702 4740 91754
rect 4684 91700 4740 91702
rect 19836 90970 19892 90972
rect 19836 90918 19838 90970
rect 19838 90918 19890 90970
rect 19890 90918 19892 90970
rect 19836 90916 19892 90918
rect 19940 90970 19996 90972
rect 19940 90918 19942 90970
rect 19942 90918 19994 90970
rect 19994 90918 19996 90970
rect 19940 90916 19996 90918
rect 20044 90970 20100 90972
rect 20044 90918 20046 90970
rect 20046 90918 20098 90970
rect 20098 90918 20100 90970
rect 20044 90916 20100 90918
rect 1820 90748 1876 90804
rect 1820 90076 1876 90132
rect 1820 82684 1876 82740
rect 1820 77362 1876 77364
rect 1820 77310 1822 77362
rect 1822 77310 1874 77362
rect 1874 77310 1876 77362
rect 1820 77308 1876 77310
rect 1820 72604 1876 72660
rect 4476 90186 4532 90188
rect 4476 90134 4478 90186
rect 4478 90134 4530 90186
rect 4530 90134 4532 90186
rect 4476 90132 4532 90134
rect 4580 90186 4636 90188
rect 4580 90134 4582 90186
rect 4582 90134 4634 90186
rect 4634 90134 4636 90186
rect 4580 90132 4636 90134
rect 4684 90186 4740 90188
rect 4684 90134 4686 90186
rect 4686 90134 4738 90186
rect 4738 90134 4740 90186
rect 4684 90132 4740 90134
rect 19836 89402 19892 89404
rect 19836 89350 19838 89402
rect 19838 89350 19890 89402
rect 19890 89350 19892 89402
rect 19836 89348 19892 89350
rect 19940 89402 19996 89404
rect 19940 89350 19942 89402
rect 19942 89350 19994 89402
rect 19994 89350 19996 89402
rect 19940 89348 19996 89350
rect 20044 89402 20100 89404
rect 20044 89350 20046 89402
rect 20046 89350 20098 89402
rect 20098 89350 20100 89402
rect 20044 89348 20100 89350
rect 4476 88618 4532 88620
rect 4476 88566 4478 88618
rect 4478 88566 4530 88618
rect 4530 88566 4532 88618
rect 4476 88564 4532 88566
rect 4580 88618 4636 88620
rect 4580 88566 4582 88618
rect 4582 88566 4634 88618
rect 4634 88566 4636 88618
rect 4580 88564 4636 88566
rect 4684 88618 4740 88620
rect 4684 88566 4686 88618
rect 4686 88566 4738 88618
rect 4738 88566 4740 88618
rect 4684 88564 4740 88566
rect 19836 87834 19892 87836
rect 19836 87782 19838 87834
rect 19838 87782 19890 87834
rect 19890 87782 19892 87834
rect 19836 87780 19892 87782
rect 19940 87834 19996 87836
rect 19940 87782 19942 87834
rect 19942 87782 19994 87834
rect 19994 87782 19996 87834
rect 19940 87780 19996 87782
rect 20044 87834 20100 87836
rect 20044 87782 20046 87834
rect 20046 87782 20098 87834
rect 20098 87782 20100 87834
rect 20044 87780 20100 87782
rect 4476 87050 4532 87052
rect 4476 86998 4478 87050
rect 4478 86998 4530 87050
rect 4530 86998 4532 87050
rect 4476 86996 4532 86998
rect 4580 87050 4636 87052
rect 4580 86998 4582 87050
rect 4582 86998 4634 87050
rect 4634 86998 4636 87050
rect 4580 86996 4636 86998
rect 4684 87050 4740 87052
rect 4684 86998 4686 87050
rect 4686 86998 4738 87050
rect 4738 86998 4740 87050
rect 4684 86996 4740 86998
rect 19836 86266 19892 86268
rect 19836 86214 19838 86266
rect 19838 86214 19890 86266
rect 19890 86214 19892 86266
rect 19836 86212 19892 86214
rect 19940 86266 19996 86268
rect 19940 86214 19942 86266
rect 19942 86214 19994 86266
rect 19994 86214 19996 86266
rect 19940 86212 19996 86214
rect 20044 86266 20100 86268
rect 20044 86214 20046 86266
rect 20046 86214 20098 86266
rect 20098 86214 20100 86266
rect 20044 86212 20100 86214
rect 4476 85482 4532 85484
rect 4476 85430 4478 85482
rect 4478 85430 4530 85482
rect 4530 85430 4532 85482
rect 4476 85428 4532 85430
rect 4580 85482 4636 85484
rect 4580 85430 4582 85482
rect 4582 85430 4634 85482
rect 4634 85430 4636 85482
rect 4580 85428 4636 85430
rect 4684 85482 4740 85484
rect 4684 85430 4686 85482
rect 4686 85430 4738 85482
rect 4738 85430 4740 85482
rect 4684 85428 4740 85430
rect 2156 84700 2212 84756
rect 2828 84812 2884 84868
rect 2492 83410 2548 83412
rect 2492 83358 2494 83410
rect 2494 83358 2546 83410
rect 2546 83358 2548 83410
rect 2492 83356 2548 83358
rect 2604 68796 2660 68852
rect 1932 67116 1988 67172
rect 1820 66556 1876 66612
rect 1820 63868 1876 63924
rect 1820 61180 1876 61236
rect 1820 57820 1876 57876
rect 3500 84866 3556 84868
rect 3500 84814 3502 84866
rect 3502 84814 3554 84866
rect 3554 84814 3556 84866
rect 3500 84812 3556 84814
rect 19836 84698 19892 84700
rect 19836 84646 19838 84698
rect 19838 84646 19890 84698
rect 19890 84646 19892 84698
rect 19836 84644 19892 84646
rect 19940 84698 19996 84700
rect 19940 84646 19942 84698
rect 19942 84646 19994 84698
rect 19994 84646 19996 84698
rect 19940 84644 19996 84646
rect 20044 84698 20100 84700
rect 20044 84646 20046 84698
rect 20046 84646 20098 84698
rect 20098 84646 20100 84698
rect 20044 84644 20100 84646
rect 4476 83914 4532 83916
rect 4476 83862 4478 83914
rect 4478 83862 4530 83914
rect 4530 83862 4532 83914
rect 4476 83860 4532 83862
rect 4580 83914 4636 83916
rect 4580 83862 4582 83914
rect 4582 83862 4634 83914
rect 4634 83862 4636 83914
rect 4580 83860 4636 83862
rect 4684 83914 4740 83916
rect 4684 83862 4686 83914
rect 4686 83862 4738 83914
rect 4738 83862 4740 83914
rect 4684 83860 4740 83862
rect 19836 83130 19892 83132
rect 19836 83078 19838 83130
rect 19838 83078 19890 83130
rect 19890 83078 19892 83130
rect 19836 83076 19892 83078
rect 19940 83130 19996 83132
rect 19940 83078 19942 83130
rect 19942 83078 19994 83130
rect 19994 83078 19996 83130
rect 19940 83076 19996 83078
rect 20044 83130 20100 83132
rect 20044 83078 20046 83130
rect 20046 83078 20098 83130
rect 20098 83078 20100 83130
rect 20044 83076 20100 83078
rect 4476 82346 4532 82348
rect 4476 82294 4478 82346
rect 4478 82294 4530 82346
rect 4530 82294 4532 82346
rect 4476 82292 4532 82294
rect 4580 82346 4636 82348
rect 4580 82294 4582 82346
rect 4582 82294 4634 82346
rect 4634 82294 4636 82346
rect 4580 82292 4636 82294
rect 4684 82346 4740 82348
rect 4684 82294 4686 82346
rect 4686 82294 4738 82346
rect 4738 82294 4740 82346
rect 4684 82292 4740 82294
rect 19836 81562 19892 81564
rect 19836 81510 19838 81562
rect 19838 81510 19890 81562
rect 19890 81510 19892 81562
rect 19836 81508 19892 81510
rect 19940 81562 19996 81564
rect 19940 81510 19942 81562
rect 19942 81510 19994 81562
rect 19994 81510 19996 81562
rect 19940 81508 19996 81510
rect 20044 81562 20100 81564
rect 20044 81510 20046 81562
rect 20046 81510 20098 81562
rect 20098 81510 20100 81562
rect 20044 81508 20100 81510
rect 4476 80778 4532 80780
rect 4476 80726 4478 80778
rect 4478 80726 4530 80778
rect 4530 80726 4532 80778
rect 4476 80724 4532 80726
rect 4580 80778 4636 80780
rect 4580 80726 4582 80778
rect 4582 80726 4634 80778
rect 4634 80726 4636 80778
rect 4580 80724 4636 80726
rect 4684 80778 4740 80780
rect 4684 80726 4686 80778
rect 4686 80726 4738 80778
rect 4738 80726 4740 80778
rect 4684 80724 4740 80726
rect 19836 79994 19892 79996
rect 19836 79942 19838 79994
rect 19838 79942 19890 79994
rect 19890 79942 19892 79994
rect 19836 79940 19892 79942
rect 19940 79994 19996 79996
rect 19940 79942 19942 79994
rect 19942 79942 19994 79994
rect 19994 79942 19996 79994
rect 19940 79940 19996 79942
rect 20044 79994 20100 79996
rect 20044 79942 20046 79994
rect 20046 79942 20098 79994
rect 20098 79942 20100 79994
rect 20044 79940 20100 79942
rect 4476 79210 4532 79212
rect 4476 79158 4478 79210
rect 4478 79158 4530 79210
rect 4530 79158 4532 79210
rect 4476 79156 4532 79158
rect 4580 79210 4636 79212
rect 4580 79158 4582 79210
rect 4582 79158 4634 79210
rect 4634 79158 4636 79210
rect 4580 79156 4636 79158
rect 4684 79210 4740 79212
rect 4684 79158 4686 79210
rect 4686 79158 4738 79210
rect 4738 79158 4740 79210
rect 4684 79156 4740 79158
rect 19836 78426 19892 78428
rect 19836 78374 19838 78426
rect 19838 78374 19890 78426
rect 19890 78374 19892 78426
rect 19836 78372 19892 78374
rect 19940 78426 19996 78428
rect 19940 78374 19942 78426
rect 19942 78374 19994 78426
rect 19994 78374 19996 78426
rect 19940 78372 19996 78374
rect 20044 78426 20100 78428
rect 20044 78374 20046 78426
rect 20046 78374 20098 78426
rect 20098 78374 20100 78426
rect 20044 78372 20100 78374
rect 4476 77642 4532 77644
rect 4476 77590 4478 77642
rect 4478 77590 4530 77642
rect 4530 77590 4532 77642
rect 4476 77588 4532 77590
rect 4580 77642 4636 77644
rect 4580 77590 4582 77642
rect 4582 77590 4634 77642
rect 4634 77590 4636 77642
rect 4580 77588 4636 77590
rect 4684 77642 4740 77644
rect 4684 77590 4686 77642
rect 4686 77590 4738 77642
rect 4738 77590 4740 77642
rect 4684 77588 4740 77590
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 3164 68850 3220 68852
rect 3164 68798 3166 68850
rect 3166 68798 3218 68850
rect 3218 68798 3220 68850
rect 3164 68796 3220 68798
rect 20076 68850 20132 68852
rect 20076 68798 20078 68850
rect 20078 68798 20130 68850
rect 20130 68798 20132 68850
rect 20076 68796 20132 68798
rect 50556 131738 50612 131740
rect 50556 131686 50558 131738
rect 50558 131686 50610 131738
rect 50610 131686 50612 131738
rect 50556 131684 50612 131686
rect 50660 131738 50716 131740
rect 50660 131686 50662 131738
rect 50662 131686 50714 131738
rect 50714 131686 50716 131738
rect 50660 131684 50716 131686
rect 50764 131738 50820 131740
rect 50764 131686 50766 131738
rect 50766 131686 50818 131738
rect 50818 131686 50820 131738
rect 50764 131684 50820 131686
rect 35196 130954 35252 130956
rect 35196 130902 35198 130954
rect 35198 130902 35250 130954
rect 35250 130902 35252 130954
rect 35196 130900 35252 130902
rect 35300 130954 35356 130956
rect 35300 130902 35302 130954
rect 35302 130902 35354 130954
rect 35354 130902 35356 130954
rect 35300 130900 35356 130902
rect 35404 130954 35460 130956
rect 35404 130902 35406 130954
rect 35406 130902 35458 130954
rect 35458 130902 35460 130954
rect 35404 130900 35460 130902
rect 50556 130170 50612 130172
rect 50556 130118 50558 130170
rect 50558 130118 50610 130170
rect 50610 130118 50612 130170
rect 50556 130116 50612 130118
rect 50660 130170 50716 130172
rect 50660 130118 50662 130170
rect 50662 130118 50714 130170
rect 50714 130118 50716 130170
rect 50660 130116 50716 130118
rect 50764 130170 50820 130172
rect 50764 130118 50766 130170
rect 50766 130118 50818 130170
rect 50818 130118 50820 130170
rect 50764 130116 50820 130118
rect 35196 129386 35252 129388
rect 35196 129334 35198 129386
rect 35198 129334 35250 129386
rect 35250 129334 35252 129386
rect 35196 129332 35252 129334
rect 35300 129386 35356 129388
rect 35300 129334 35302 129386
rect 35302 129334 35354 129386
rect 35354 129334 35356 129386
rect 35300 129332 35356 129334
rect 35404 129386 35460 129388
rect 35404 129334 35406 129386
rect 35406 129334 35458 129386
rect 35458 129334 35460 129386
rect 35404 129332 35460 129334
rect 50556 128602 50612 128604
rect 50556 128550 50558 128602
rect 50558 128550 50610 128602
rect 50610 128550 50612 128602
rect 50556 128548 50612 128550
rect 50660 128602 50716 128604
rect 50660 128550 50662 128602
rect 50662 128550 50714 128602
rect 50714 128550 50716 128602
rect 50660 128548 50716 128550
rect 50764 128602 50820 128604
rect 50764 128550 50766 128602
rect 50766 128550 50818 128602
rect 50818 128550 50820 128602
rect 50764 128548 50820 128550
rect 35196 127818 35252 127820
rect 35196 127766 35198 127818
rect 35198 127766 35250 127818
rect 35250 127766 35252 127818
rect 35196 127764 35252 127766
rect 35300 127818 35356 127820
rect 35300 127766 35302 127818
rect 35302 127766 35354 127818
rect 35354 127766 35356 127818
rect 35300 127764 35356 127766
rect 35404 127818 35460 127820
rect 35404 127766 35406 127818
rect 35406 127766 35458 127818
rect 35458 127766 35460 127818
rect 35404 127764 35460 127766
rect 50556 127034 50612 127036
rect 50556 126982 50558 127034
rect 50558 126982 50610 127034
rect 50610 126982 50612 127034
rect 50556 126980 50612 126982
rect 50660 127034 50716 127036
rect 50660 126982 50662 127034
rect 50662 126982 50714 127034
rect 50714 126982 50716 127034
rect 50660 126980 50716 126982
rect 50764 127034 50820 127036
rect 50764 126982 50766 127034
rect 50766 126982 50818 127034
rect 50818 126982 50820 127034
rect 50764 126980 50820 126982
rect 35196 126250 35252 126252
rect 35196 126198 35198 126250
rect 35198 126198 35250 126250
rect 35250 126198 35252 126250
rect 35196 126196 35252 126198
rect 35300 126250 35356 126252
rect 35300 126198 35302 126250
rect 35302 126198 35354 126250
rect 35354 126198 35356 126250
rect 35300 126196 35356 126198
rect 35404 126250 35460 126252
rect 35404 126198 35406 126250
rect 35406 126198 35458 126250
rect 35458 126198 35460 126250
rect 35404 126196 35460 126198
rect 50556 125466 50612 125468
rect 50556 125414 50558 125466
rect 50558 125414 50610 125466
rect 50610 125414 50612 125466
rect 50556 125412 50612 125414
rect 50660 125466 50716 125468
rect 50660 125414 50662 125466
rect 50662 125414 50714 125466
rect 50714 125414 50716 125466
rect 50660 125412 50716 125414
rect 50764 125466 50820 125468
rect 50764 125414 50766 125466
rect 50766 125414 50818 125466
rect 50818 125414 50820 125466
rect 50764 125412 50820 125414
rect 35196 124682 35252 124684
rect 35196 124630 35198 124682
rect 35198 124630 35250 124682
rect 35250 124630 35252 124682
rect 35196 124628 35252 124630
rect 35300 124682 35356 124684
rect 35300 124630 35302 124682
rect 35302 124630 35354 124682
rect 35354 124630 35356 124682
rect 35300 124628 35356 124630
rect 35404 124682 35460 124684
rect 35404 124630 35406 124682
rect 35406 124630 35458 124682
rect 35458 124630 35460 124682
rect 35404 124628 35460 124630
rect 50556 123898 50612 123900
rect 50556 123846 50558 123898
rect 50558 123846 50610 123898
rect 50610 123846 50612 123898
rect 50556 123844 50612 123846
rect 50660 123898 50716 123900
rect 50660 123846 50662 123898
rect 50662 123846 50714 123898
rect 50714 123846 50716 123898
rect 50660 123844 50716 123846
rect 50764 123898 50820 123900
rect 50764 123846 50766 123898
rect 50766 123846 50818 123898
rect 50818 123846 50820 123898
rect 50764 123844 50820 123846
rect 35196 123114 35252 123116
rect 35196 123062 35198 123114
rect 35198 123062 35250 123114
rect 35250 123062 35252 123114
rect 35196 123060 35252 123062
rect 35300 123114 35356 123116
rect 35300 123062 35302 123114
rect 35302 123062 35354 123114
rect 35354 123062 35356 123114
rect 35300 123060 35356 123062
rect 35404 123114 35460 123116
rect 35404 123062 35406 123114
rect 35406 123062 35458 123114
rect 35458 123062 35460 123114
rect 35404 123060 35460 123062
rect 50556 122330 50612 122332
rect 50556 122278 50558 122330
rect 50558 122278 50610 122330
rect 50610 122278 50612 122330
rect 50556 122276 50612 122278
rect 50660 122330 50716 122332
rect 50660 122278 50662 122330
rect 50662 122278 50714 122330
rect 50714 122278 50716 122330
rect 50660 122276 50716 122278
rect 50764 122330 50820 122332
rect 50764 122278 50766 122330
rect 50766 122278 50818 122330
rect 50818 122278 50820 122330
rect 50764 122276 50820 122278
rect 35196 121546 35252 121548
rect 35196 121494 35198 121546
rect 35198 121494 35250 121546
rect 35250 121494 35252 121546
rect 35196 121492 35252 121494
rect 35300 121546 35356 121548
rect 35300 121494 35302 121546
rect 35302 121494 35354 121546
rect 35354 121494 35356 121546
rect 35300 121492 35356 121494
rect 35404 121546 35460 121548
rect 35404 121494 35406 121546
rect 35406 121494 35458 121546
rect 35458 121494 35460 121546
rect 35404 121492 35460 121494
rect 50556 120762 50612 120764
rect 50556 120710 50558 120762
rect 50558 120710 50610 120762
rect 50610 120710 50612 120762
rect 50556 120708 50612 120710
rect 50660 120762 50716 120764
rect 50660 120710 50662 120762
rect 50662 120710 50714 120762
rect 50714 120710 50716 120762
rect 50660 120708 50716 120710
rect 50764 120762 50820 120764
rect 50764 120710 50766 120762
rect 50766 120710 50818 120762
rect 50818 120710 50820 120762
rect 50764 120708 50820 120710
rect 35196 119978 35252 119980
rect 35196 119926 35198 119978
rect 35198 119926 35250 119978
rect 35250 119926 35252 119978
rect 35196 119924 35252 119926
rect 35300 119978 35356 119980
rect 35300 119926 35302 119978
rect 35302 119926 35354 119978
rect 35354 119926 35356 119978
rect 35300 119924 35356 119926
rect 35404 119978 35460 119980
rect 35404 119926 35406 119978
rect 35406 119926 35458 119978
rect 35458 119926 35460 119978
rect 35404 119924 35460 119926
rect 50556 119194 50612 119196
rect 50556 119142 50558 119194
rect 50558 119142 50610 119194
rect 50610 119142 50612 119194
rect 50556 119140 50612 119142
rect 50660 119194 50716 119196
rect 50660 119142 50662 119194
rect 50662 119142 50714 119194
rect 50714 119142 50716 119194
rect 50660 119140 50716 119142
rect 50764 119194 50820 119196
rect 50764 119142 50766 119194
rect 50766 119142 50818 119194
rect 50818 119142 50820 119194
rect 50764 119140 50820 119142
rect 35196 118410 35252 118412
rect 35196 118358 35198 118410
rect 35198 118358 35250 118410
rect 35250 118358 35252 118410
rect 35196 118356 35252 118358
rect 35300 118410 35356 118412
rect 35300 118358 35302 118410
rect 35302 118358 35354 118410
rect 35354 118358 35356 118410
rect 35300 118356 35356 118358
rect 35404 118410 35460 118412
rect 35404 118358 35406 118410
rect 35406 118358 35458 118410
rect 35458 118358 35460 118410
rect 35404 118356 35460 118358
rect 50556 117626 50612 117628
rect 50556 117574 50558 117626
rect 50558 117574 50610 117626
rect 50610 117574 50612 117626
rect 50556 117572 50612 117574
rect 50660 117626 50716 117628
rect 50660 117574 50662 117626
rect 50662 117574 50714 117626
rect 50714 117574 50716 117626
rect 50660 117572 50716 117574
rect 50764 117626 50820 117628
rect 50764 117574 50766 117626
rect 50766 117574 50818 117626
rect 50818 117574 50820 117626
rect 50764 117572 50820 117574
rect 35196 116842 35252 116844
rect 35196 116790 35198 116842
rect 35198 116790 35250 116842
rect 35250 116790 35252 116842
rect 35196 116788 35252 116790
rect 35300 116842 35356 116844
rect 35300 116790 35302 116842
rect 35302 116790 35354 116842
rect 35354 116790 35356 116842
rect 35300 116788 35356 116790
rect 35404 116842 35460 116844
rect 35404 116790 35406 116842
rect 35406 116790 35458 116842
rect 35458 116790 35460 116842
rect 35404 116788 35460 116790
rect 50556 116058 50612 116060
rect 50556 116006 50558 116058
rect 50558 116006 50610 116058
rect 50610 116006 50612 116058
rect 50556 116004 50612 116006
rect 50660 116058 50716 116060
rect 50660 116006 50662 116058
rect 50662 116006 50714 116058
rect 50714 116006 50716 116058
rect 50660 116004 50716 116006
rect 50764 116058 50820 116060
rect 50764 116006 50766 116058
rect 50766 116006 50818 116058
rect 50818 116006 50820 116058
rect 50764 116004 50820 116006
rect 35196 115274 35252 115276
rect 35196 115222 35198 115274
rect 35198 115222 35250 115274
rect 35250 115222 35252 115274
rect 35196 115220 35252 115222
rect 35300 115274 35356 115276
rect 35300 115222 35302 115274
rect 35302 115222 35354 115274
rect 35354 115222 35356 115274
rect 35300 115220 35356 115222
rect 35404 115274 35460 115276
rect 35404 115222 35406 115274
rect 35406 115222 35458 115274
rect 35458 115222 35460 115274
rect 35404 115220 35460 115222
rect 50556 114490 50612 114492
rect 50556 114438 50558 114490
rect 50558 114438 50610 114490
rect 50610 114438 50612 114490
rect 50556 114436 50612 114438
rect 50660 114490 50716 114492
rect 50660 114438 50662 114490
rect 50662 114438 50714 114490
rect 50714 114438 50716 114490
rect 50660 114436 50716 114438
rect 50764 114490 50820 114492
rect 50764 114438 50766 114490
rect 50766 114438 50818 114490
rect 50818 114438 50820 114490
rect 50764 114436 50820 114438
rect 35196 113706 35252 113708
rect 35196 113654 35198 113706
rect 35198 113654 35250 113706
rect 35250 113654 35252 113706
rect 35196 113652 35252 113654
rect 35300 113706 35356 113708
rect 35300 113654 35302 113706
rect 35302 113654 35354 113706
rect 35354 113654 35356 113706
rect 35300 113652 35356 113654
rect 35404 113706 35460 113708
rect 35404 113654 35406 113706
rect 35406 113654 35458 113706
rect 35458 113654 35460 113706
rect 35404 113652 35460 113654
rect 50556 112922 50612 112924
rect 50556 112870 50558 112922
rect 50558 112870 50610 112922
rect 50610 112870 50612 112922
rect 50556 112868 50612 112870
rect 50660 112922 50716 112924
rect 50660 112870 50662 112922
rect 50662 112870 50714 112922
rect 50714 112870 50716 112922
rect 50660 112868 50716 112870
rect 50764 112922 50820 112924
rect 50764 112870 50766 112922
rect 50766 112870 50818 112922
rect 50818 112870 50820 112922
rect 50764 112868 50820 112870
rect 35196 112138 35252 112140
rect 35196 112086 35198 112138
rect 35198 112086 35250 112138
rect 35250 112086 35252 112138
rect 35196 112084 35252 112086
rect 35300 112138 35356 112140
rect 35300 112086 35302 112138
rect 35302 112086 35354 112138
rect 35354 112086 35356 112138
rect 35300 112084 35356 112086
rect 35404 112138 35460 112140
rect 35404 112086 35406 112138
rect 35406 112086 35458 112138
rect 35458 112086 35460 112138
rect 35404 112084 35460 112086
rect 50556 111354 50612 111356
rect 50556 111302 50558 111354
rect 50558 111302 50610 111354
rect 50610 111302 50612 111354
rect 50556 111300 50612 111302
rect 50660 111354 50716 111356
rect 50660 111302 50662 111354
rect 50662 111302 50714 111354
rect 50714 111302 50716 111354
rect 50660 111300 50716 111302
rect 50764 111354 50820 111356
rect 50764 111302 50766 111354
rect 50766 111302 50818 111354
rect 50818 111302 50820 111354
rect 50764 111300 50820 111302
rect 35196 110570 35252 110572
rect 35196 110518 35198 110570
rect 35198 110518 35250 110570
rect 35250 110518 35252 110570
rect 35196 110516 35252 110518
rect 35300 110570 35356 110572
rect 35300 110518 35302 110570
rect 35302 110518 35354 110570
rect 35354 110518 35356 110570
rect 35300 110516 35356 110518
rect 35404 110570 35460 110572
rect 35404 110518 35406 110570
rect 35406 110518 35458 110570
rect 35458 110518 35460 110570
rect 35404 110516 35460 110518
rect 50556 109786 50612 109788
rect 50556 109734 50558 109786
rect 50558 109734 50610 109786
rect 50610 109734 50612 109786
rect 50556 109732 50612 109734
rect 50660 109786 50716 109788
rect 50660 109734 50662 109786
rect 50662 109734 50714 109786
rect 50714 109734 50716 109786
rect 50660 109732 50716 109734
rect 50764 109786 50820 109788
rect 50764 109734 50766 109786
rect 50766 109734 50818 109786
rect 50818 109734 50820 109786
rect 50764 109732 50820 109734
rect 35196 109002 35252 109004
rect 35196 108950 35198 109002
rect 35198 108950 35250 109002
rect 35250 108950 35252 109002
rect 35196 108948 35252 108950
rect 35300 109002 35356 109004
rect 35300 108950 35302 109002
rect 35302 108950 35354 109002
rect 35354 108950 35356 109002
rect 35300 108948 35356 108950
rect 35404 109002 35460 109004
rect 35404 108950 35406 109002
rect 35406 108950 35458 109002
rect 35458 108950 35460 109002
rect 35404 108948 35460 108950
rect 50556 108218 50612 108220
rect 50556 108166 50558 108218
rect 50558 108166 50610 108218
rect 50610 108166 50612 108218
rect 50556 108164 50612 108166
rect 50660 108218 50716 108220
rect 50660 108166 50662 108218
rect 50662 108166 50714 108218
rect 50714 108166 50716 108218
rect 50660 108164 50716 108166
rect 50764 108218 50820 108220
rect 50764 108166 50766 108218
rect 50766 108166 50818 108218
rect 50818 108166 50820 108218
rect 50764 108164 50820 108166
rect 35196 107434 35252 107436
rect 35196 107382 35198 107434
rect 35198 107382 35250 107434
rect 35250 107382 35252 107434
rect 35196 107380 35252 107382
rect 35300 107434 35356 107436
rect 35300 107382 35302 107434
rect 35302 107382 35354 107434
rect 35354 107382 35356 107434
rect 35300 107380 35356 107382
rect 35404 107434 35460 107436
rect 35404 107382 35406 107434
rect 35406 107382 35458 107434
rect 35458 107382 35460 107434
rect 35404 107380 35460 107382
rect 50556 106650 50612 106652
rect 50556 106598 50558 106650
rect 50558 106598 50610 106650
rect 50610 106598 50612 106650
rect 50556 106596 50612 106598
rect 50660 106650 50716 106652
rect 50660 106598 50662 106650
rect 50662 106598 50714 106650
rect 50714 106598 50716 106650
rect 50660 106596 50716 106598
rect 50764 106650 50820 106652
rect 50764 106598 50766 106650
rect 50766 106598 50818 106650
rect 50818 106598 50820 106650
rect 50764 106596 50820 106598
rect 35196 105866 35252 105868
rect 35196 105814 35198 105866
rect 35198 105814 35250 105866
rect 35250 105814 35252 105866
rect 35196 105812 35252 105814
rect 35300 105866 35356 105868
rect 35300 105814 35302 105866
rect 35302 105814 35354 105866
rect 35354 105814 35356 105866
rect 35300 105812 35356 105814
rect 35404 105866 35460 105868
rect 35404 105814 35406 105866
rect 35406 105814 35458 105866
rect 35458 105814 35460 105866
rect 35404 105812 35460 105814
rect 50556 105082 50612 105084
rect 50556 105030 50558 105082
rect 50558 105030 50610 105082
rect 50610 105030 50612 105082
rect 50556 105028 50612 105030
rect 50660 105082 50716 105084
rect 50660 105030 50662 105082
rect 50662 105030 50714 105082
rect 50714 105030 50716 105082
rect 50660 105028 50716 105030
rect 50764 105082 50820 105084
rect 50764 105030 50766 105082
rect 50766 105030 50818 105082
rect 50818 105030 50820 105082
rect 50764 105028 50820 105030
rect 35196 104298 35252 104300
rect 35196 104246 35198 104298
rect 35198 104246 35250 104298
rect 35250 104246 35252 104298
rect 35196 104244 35252 104246
rect 35300 104298 35356 104300
rect 35300 104246 35302 104298
rect 35302 104246 35354 104298
rect 35354 104246 35356 104298
rect 35300 104244 35356 104246
rect 35404 104298 35460 104300
rect 35404 104246 35406 104298
rect 35406 104246 35458 104298
rect 35458 104246 35460 104298
rect 35404 104244 35460 104246
rect 50556 103514 50612 103516
rect 50556 103462 50558 103514
rect 50558 103462 50610 103514
rect 50610 103462 50612 103514
rect 50556 103460 50612 103462
rect 50660 103514 50716 103516
rect 50660 103462 50662 103514
rect 50662 103462 50714 103514
rect 50714 103462 50716 103514
rect 50660 103460 50716 103462
rect 50764 103514 50820 103516
rect 50764 103462 50766 103514
rect 50766 103462 50818 103514
rect 50818 103462 50820 103514
rect 50764 103460 50820 103462
rect 35196 102730 35252 102732
rect 35196 102678 35198 102730
rect 35198 102678 35250 102730
rect 35250 102678 35252 102730
rect 35196 102676 35252 102678
rect 35300 102730 35356 102732
rect 35300 102678 35302 102730
rect 35302 102678 35354 102730
rect 35354 102678 35356 102730
rect 35300 102676 35356 102678
rect 35404 102730 35460 102732
rect 35404 102678 35406 102730
rect 35406 102678 35458 102730
rect 35458 102678 35460 102730
rect 35404 102676 35460 102678
rect 50556 101946 50612 101948
rect 50556 101894 50558 101946
rect 50558 101894 50610 101946
rect 50610 101894 50612 101946
rect 50556 101892 50612 101894
rect 50660 101946 50716 101948
rect 50660 101894 50662 101946
rect 50662 101894 50714 101946
rect 50714 101894 50716 101946
rect 50660 101892 50716 101894
rect 50764 101946 50820 101948
rect 50764 101894 50766 101946
rect 50766 101894 50818 101946
rect 50818 101894 50820 101946
rect 50764 101892 50820 101894
rect 35196 101162 35252 101164
rect 35196 101110 35198 101162
rect 35198 101110 35250 101162
rect 35250 101110 35252 101162
rect 35196 101108 35252 101110
rect 35300 101162 35356 101164
rect 35300 101110 35302 101162
rect 35302 101110 35354 101162
rect 35354 101110 35356 101162
rect 35300 101108 35356 101110
rect 35404 101162 35460 101164
rect 35404 101110 35406 101162
rect 35406 101110 35458 101162
rect 35458 101110 35460 101162
rect 35404 101108 35460 101110
rect 50556 100378 50612 100380
rect 50556 100326 50558 100378
rect 50558 100326 50610 100378
rect 50610 100326 50612 100378
rect 50556 100324 50612 100326
rect 50660 100378 50716 100380
rect 50660 100326 50662 100378
rect 50662 100326 50714 100378
rect 50714 100326 50716 100378
rect 50660 100324 50716 100326
rect 50764 100378 50820 100380
rect 50764 100326 50766 100378
rect 50766 100326 50818 100378
rect 50818 100326 50820 100378
rect 50764 100324 50820 100326
rect 35196 99594 35252 99596
rect 35196 99542 35198 99594
rect 35198 99542 35250 99594
rect 35250 99542 35252 99594
rect 35196 99540 35252 99542
rect 35300 99594 35356 99596
rect 35300 99542 35302 99594
rect 35302 99542 35354 99594
rect 35354 99542 35356 99594
rect 35300 99540 35356 99542
rect 35404 99594 35460 99596
rect 35404 99542 35406 99594
rect 35406 99542 35458 99594
rect 35458 99542 35460 99594
rect 35404 99540 35460 99542
rect 50556 98810 50612 98812
rect 50556 98758 50558 98810
rect 50558 98758 50610 98810
rect 50610 98758 50612 98810
rect 50556 98756 50612 98758
rect 50660 98810 50716 98812
rect 50660 98758 50662 98810
rect 50662 98758 50714 98810
rect 50714 98758 50716 98810
rect 50660 98756 50716 98758
rect 50764 98810 50820 98812
rect 50764 98758 50766 98810
rect 50766 98758 50818 98810
rect 50818 98758 50820 98810
rect 50764 98756 50820 98758
rect 35196 98026 35252 98028
rect 35196 97974 35198 98026
rect 35198 97974 35250 98026
rect 35250 97974 35252 98026
rect 35196 97972 35252 97974
rect 35300 98026 35356 98028
rect 35300 97974 35302 98026
rect 35302 97974 35354 98026
rect 35354 97974 35356 98026
rect 35300 97972 35356 97974
rect 35404 98026 35460 98028
rect 35404 97974 35406 98026
rect 35406 97974 35458 98026
rect 35458 97974 35460 98026
rect 35404 97972 35460 97974
rect 50556 97242 50612 97244
rect 50556 97190 50558 97242
rect 50558 97190 50610 97242
rect 50610 97190 50612 97242
rect 50556 97188 50612 97190
rect 50660 97242 50716 97244
rect 50660 97190 50662 97242
rect 50662 97190 50714 97242
rect 50714 97190 50716 97242
rect 50660 97188 50716 97190
rect 50764 97242 50820 97244
rect 50764 97190 50766 97242
rect 50766 97190 50818 97242
rect 50818 97190 50820 97242
rect 50764 97188 50820 97190
rect 35196 96458 35252 96460
rect 35196 96406 35198 96458
rect 35198 96406 35250 96458
rect 35250 96406 35252 96458
rect 35196 96404 35252 96406
rect 35300 96458 35356 96460
rect 35300 96406 35302 96458
rect 35302 96406 35354 96458
rect 35354 96406 35356 96458
rect 35300 96404 35356 96406
rect 35404 96458 35460 96460
rect 35404 96406 35406 96458
rect 35406 96406 35458 96458
rect 35458 96406 35460 96458
rect 35404 96404 35460 96406
rect 50556 95674 50612 95676
rect 50556 95622 50558 95674
rect 50558 95622 50610 95674
rect 50610 95622 50612 95674
rect 50556 95620 50612 95622
rect 50660 95674 50716 95676
rect 50660 95622 50662 95674
rect 50662 95622 50714 95674
rect 50714 95622 50716 95674
rect 50660 95620 50716 95622
rect 50764 95674 50820 95676
rect 50764 95622 50766 95674
rect 50766 95622 50818 95674
rect 50818 95622 50820 95674
rect 50764 95620 50820 95622
rect 35196 94890 35252 94892
rect 35196 94838 35198 94890
rect 35198 94838 35250 94890
rect 35250 94838 35252 94890
rect 35196 94836 35252 94838
rect 35300 94890 35356 94892
rect 35300 94838 35302 94890
rect 35302 94838 35354 94890
rect 35354 94838 35356 94890
rect 35300 94836 35356 94838
rect 35404 94890 35460 94892
rect 35404 94838 35406 94890
rect 35406 94838 35458 94890
rect 35458 94838 35460 94890
rect 35404 94836 35460 94838
rect 50556 94106 50612 94108
rect 50556 94054 50558 94106
rect 50558 94054 50610 94106
rect 50610 94054 50612 94106
rect 50556 94052 50612 94054
rect 50660 94106 50716 94108
rect 50660 94054 50662 94106
rect 50662 94054 50714 94106
rect 50714 94054 50716 94106
rect 50660 94052 50716 94054
rect 50764 94106 50820 94108
rect 50764 94054 50766 94106
rect 50766 94054 50818 94106
rect 50818 94054 50820 94106
rect 50764 94052 50820 94054
rect 35196 93322 35252 93324
rect 35196 93270 35198 93322
rect 35198 93270 35250 93322
rect 35250 93270 35252 93322
rect 35196 93268 35252 93270
rect 35300 93322 35356 93324
rect 35300 93270 35302 93322
rect 35302 93270 35354 93322
rect 35354 93270 35356 93322
rect 35300 93268 35356 93270
rect 35404 93322 35460 93324
rect 35404 93270 35406 93322
rect 35406 93270 35458 93322
rect 35458 93270 35460 93322
rect 35404 93268 35460 93270
rect 50556 92538 50612 92540
rect 50556 92486 50558 92538
rect 50558 92486 50610 92538
rect 50610 92486 50612 92538
rect 50556 92484 50612 92486
rect 50660 92538 50716 92540
rect 50660 92486 50662 92538
rect 50662 92486 50714 92538
rect 50714 92486 50716 92538
rect 50660 92484 50716 92486
rect 50764 92538 50820 92540
rect 50764 92486 50766 92538
rect 50766 92486 50818 92538
rect 50818 92486 50820 92538
rect 50764 92484 50820 92486
rect 35196 91754 35252 91756
rect 35196 91702 35198 91754
rect 35198 91702 35250 91754
rect 35250 91702 35252 91754
rect 35196 91700 35252 91702
rect 35300 91754 35356 91756
rect 35300 91702 35302 91754
rect 35302 91702 35354 91754
rect 35354 91702 35356 91754
rect 35300 91700 35356 91702
rect 35404 91754 35460 91756
rect 35404 91702 35406 91754
rect 35406 91702 35458 91754
rect 35458 91702 35460 91754
rect 35404 91700 35460 91702
rect 50556 90970 50612 90972
rect 50556 90918 50558 90970
rect 50558 90918 50610 90970
rect 50610 90918 50612 90970
rect 50556 90916 50612 90918
rect 50660 90970 50716 90972
rect 50660 90918 50662 90970
rect 50662 90918 50714 90970
rect 50714 90918 50716 90970
rect 50660 90916 50716 90918
rect 50764 90970 50820 90972
rect 50764 90918 50766 90970
rect 50766 90918 50818 90970
rect 50818 90918 50820 90970
rect 50764 90916 50820 90918
rect 35196 90186 35252 90188
rect 35196 90134 35198 90186
rect 35198 90134 35250 90186
rect 35250 90134 35252 90186
rect 35196 90132 35252 90134
rect 35300 90186 35356 90188
rect 35300 90134 35302 90186
rect 35302 90134 35354 90186
rect 35354 90134 35356 90186
rect 35300 90132 35356 90134
rect 35404 90186 35460 90188
rect 35404 90134 35406 90186
rect 35406 90134 35458 90186
rect 35458 90134 35460 90186
rect 35404 90132 35460 90134
rect 50556 89402 50612 89404
rect 50556 89350 50558 89402
rect 50558 89350 50610 89402
rect 50610 89350 50612 89402
rect 50556 89348 50612 89350
rect 50660 89402 50716 89404
rect 50660 89350 50662 89402
rect 50662 89350 50714 89402
rect 50714 89350 50716 89402
rect 50660 89348 50716 89350
rect 50764 89402 50820 89404
rect 50764 89350 50766 89402
rect 50766 89350 50818 89402
rect 50818 89350 50820 89402
rect 50764 89348 50820 89350
rect 35196 88618 35252 88620
rect 35196 88566 35198 88618
rect 35198 88566 35250 88618
rect 35250 88566 35252 88618
rect 35196 88564 35252 88566
rect 35300 88618 35356 88620
rect 35300 88566 35302 88618
rect 35302 88566 35354 88618
rect 35354 88566 35356 88618
rect 35300 88564 35356 88566
rect 35404 88618 35460 88620
rect 35404 88566 35406 88618
rect 35406 88566 35458 88618
rect 35458 88566 35460 88618
rect 35404 88564 35460 88566
rect 50556 87834 50612 87836
rect 50556 87782 50558 87834
rect 50558 87782 50610 87834
rect 50610 87782 50612 87834
rect 50556 87780 50612 87782
rect 50660 87834 50716 87836
rect 50660 87782 50662 87834
rect 50662 87782 50714 87834
rect 50714 87782 50716 87834
rect 50660 87780 50716 87782
rect 50764 87834 50820 87836
rect 50764 87782 50766 87834
rect 50766 87782 50818 87834
rect 50818 87782 50820 87834
rect 50764 87780 50820 87782
rect 35196 87050 35252 87052
rect 35196 86998 35198 87050
rect 35198 86998 35250 87050
rect 35250 86998 35252 87050
rect 35196 86996 35252 86998
rect 35300 87050 35356 87052
rect 35300 86998 35302 87050
rect 35302 86998 35354 87050
rect 35354 86998 35356 87050
rect 35300 86996 35356 86998
rect 35404 87050 35460 87052
rect 35404 86998 35406 87050
rect 35406 86998 35458 87050
rect 35458 86998 35460 87050
rect 35404 86996 35460 86998
rect 50556 86266 50612 86268
rect 50556 86214 50558 86266
rect 50558 86214 50610 86266
rect 50610 86214 50612 86266
rect 50556 86212 50612 86214
rect 50660 86266 50716 86268
rect 50660 86214 50662 86266
rect 50662 86214 50714 86266
rect 50714 86214 50716 86266
rect 50660 86212 50716 86214
rect 50764 86266 50820 86268
rect 50764 86214 50766 86266
rect 50766 86214 50818 86266
rect 50818 86214 50820 86266
rect 50764 86212 50820 86214
rect 35196 85482 35252 85484
rect 35196 85430 35198 85482
rect 35198 85430 35250 85482
rect 35250 85430 35252 85482
rect 35196 85428 35252 85430
rect 35300 85482 35356 85484
rect 35300 85430 35302 85482
rect 35302 85430 35354 85482
rect 35354 85430 35356 85482
rect 35300 85428 35356 85430
rect 35404 85482 35460 85484
rect 35404 85430 35406 85482
rect 35406 85430 35458 85482
rect 35458 85430 35460 85482
rect 35404 85428 35460 85430
rect 50556 84698 50612 84700
rect 50556 84646 50558 84698
rect 50558 84646 50610 84698
rect 50610 84646 50612 84698
rect 50556 84644 50612 84646
rect 50660 84698 50716 84700
rect 50660 84646 50662 84698
rect 50662 84646 50714 84698
rect 50714 84646 50716 84698
rect 50660 84644 50716 84646
rect 50764 84698 50820 84700
rect 50764 84646 50766 84698
rect 50766 84646 50818 84698
rect 50818 84646 50820 84698
rect 50764 84644 50820 84646
rect 35196 83914 35252 83916
rect 35196 83862 35198 83914
rect 35198 83862 35250 83914
rect 35250 83862 35252 83914
rect 35196 83860 35252 83862
rect 35300 83914 35356 83916
rect 35300 83862 35302 83914
rect 35302 83862 35354 83914
rect 35354 83862 35356 83914
rect 35300 83860 35356 83862
rect 35404 83914 35460 83916
rect 35404 83862 35406 83914
rect 35406 83862 35458 83914
rect 35458 83862 35460 83914
rect 35404 83860 35460 83862
rect 50556 83130 50612 83132
rect 50556 83078 50558 83130
rect 50558 83078 50610 83130
rect 50610 83078 50612 83130
rect 50556 83076 50612 83078
rect 50660 83130 50716 83132
rect 50660 83078 50662 83130
rect 50662 83078 50714 83130
rect 50714 83078 50716 83130
rect 50660 83076 50716 83078
rect 50764 83130 50820 83132
rect 50764 83078 50766 83130
rect 50766 83078 50818 83130
rect 50818 83078 50820 83130
rect 50764 83076 50820 83078
rect 35196 82346 35252 82348
rect 35196 82294 35198 82346
rect 35198 82294 35250 82346
rect 35250 82294 35252 82346
rect 35196 82292 35252 82294
rect 35300 82346 35356 82348
rect 35300 82294 35302 82346
rect 35302 82294 35354 82346
rect 35354 82294 35356 82346
rect 35300 82292 35356 82294
rect 35404 82346 35460 82348
rect 35404 82294 35406 82346
rect 35406 82294 35458 82346
rect 35458 82294 35460 82346
rect 35404 82292 35460 82294
rect 50556 81562 50612 81564
rect 50556 81510 50558 81562
rect 50558 81510 50610 81562
rect 50610 81510 50612 81562
rect 50556 81508 50612 81510
rect 50660 81562 50716 81564
rect 50660 81510 50662 81562
rect 50662 81510 50714 81562
rect 50714 81510 50716 81562
rect 50660 81508 50716 81510
rect 50764 81562 50820 81564
rect 50764 81510 50766 81562
rect 50766 81510 50818 81562
rect 50818 81510 50820 81562
rect 50764 81508 50820 81510
rect 35196 80778 35252 80780
rect 35196 80726 35198 80778
rect 35198 80726 35250 80778
rect 35250 80726 35252 80778
rect 35196 80724 35252 80726
rect 35300 80778 35356 80780
rect 35300 80726 35302 80778
rect 35302 80726 35354 80778
rect 35354 80726 35356 80778
rect 35300 80724 35356 80726
rect 35404 80778 35460 80780
rect 35404 80726 35406 80778
rect 35406 80726 35458 80778
rect 35458 80726 35460 80778
rect 35404 80724 35460 80726
rect 50556 79994 50612 79996
rect 50556 79942 50558 79994
rect 50558 79942 50610 79994
rect 50610 79942 50612 79994
rect 50556 79940 50612 79942
rect 50660 79994 50716 79996
rect 50660 79942 50662 79994
rect 50662 79942 50714 79994
rect 50714 79942 50716 79994
rect 50660 79940 50716 79942
rect 50764 79994 50820 79996
rect 50764 79942 50766 79994
rect 50766 79942 50818 79994
rect 50818 79942 50820 79994
rect 50764 79940 50820 79942
rect 35196 79210 35252 79212
rect 35196 79158 35198 79210
rect 35198 79158 35250 79210
rect 35250 79158 35252 79210
rect 35196 79156 35252 79158
rect 35300 79210 35356 79212
rect 35300 79158 35302 79210
rect 35302 79158 35354 79210
rect 35354 79158 35356 79210
rect 35300 79156 35356 79158
rect 35404 79210 35460 79212
rect 35404 79158 35406 79210
rect 35406 79158 35458 79210
rect 35458 79158 35460 79210
rect 35404 79156 35460 79158
rect 50556 78426 50612 78428
rect 50556 78374 50558 78426
rect 50558 78374 50610 78426
rect 50610 78374 50612 78426
rect 50556 78372 50612 78374
rect 50660 78426 50716 78428
rect 50660 78374 50662 78426
rect 50662 78374 50714 78426
rect 50714 78374 50716 78426
rect 50660 78372 50716 78374
rect 50764 78426 50820 78428
rect 50764 78374 50766 78426
rect 50766 78374 50818 78426
rect 50818 78374 50820 78426
rect 50764 78372 50820 78374
rect 35196 77642 35252 77644
rect 35196 77590 35198 77642
rect 35198 77590 35250 77642
rect 35250 77590 35252 77642
rect 35196 77588 35252 77590
rect 35300 77642 35356 77644
rect 35300 77590 35302 77642
rect 35302 77590 35354 77642
rect 35354 77590 35356 77642
rect 35300 77588 35356 77590
rect 35404 77642 35460 77644
rect 35404 77590 35406 77642
rect 35406 77590 35458 77642
rect 35458 77590 35460 77642
rect 35404 77588 35460 77590
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 21420 68796 21476 68852
rect 19964 68514 20020 68516
rect 19964 68462 19966 68514
rect 19966 68462 20018 68514
rect 20018 68462 20020 68514
rect 19964 68460 20020 68462
rect 20636 68514 20692 68516
rect 20636 68462 20638 68514
rect 20638 68462 20690 68514
rect 20690 68462 20692 68514
rect 20636 68460 20692 68462
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 2716 67564 2772 67620
rect 3500 67618 3556 67620
rect 3500 67566 3502 67618
rect 3502 67566 3554 67618
rect 3554 67566 3556 67618
rect 3500 67564 3556 67566
rect 3724 67004 3780 67060
rect 1820 52444 1876 52500
rect 1820 49084 1876 49140
rect 3052 48076 3108 48132
rect 3500 48130 3556 48132
rect 3500 48078 3502 48130
rect 3502 48078 3554 48130
rect 3554 48078 3556 48130
rect 3500 48076 3556 48078
rect 2044 47740 2100 47796
rect 1820 46396 1876 46452
rect 2156 45330 2212 45332
rect 2156 45278 2158 45330
rect 2158 45278 2210 45330
rect 2210 45278 2212 45330
rect 2156 45276 2212 45278
rect 1932 45052 1988 45108
rect 1820 44434 1876 44436
rect 1820 44382 1822 44434
rect 1822 44382 1874 44434
rect 1874 44382 1876 44434
rect 1820 44380 1876 44382
rect 1820 41692 1876 41748
rect 5068 67564 5124 67620
rect 4620 67058 4676 67060
rect 4620 67006 4622 67058
rect 4622 67006 4674 67058
rect 4674 67006 4676 67058
rect 4620 67004 4676 67006
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 6300 67170 6356 67172
rect 6300 67118 6302 67170
rect 6302 67118 6354 67170
rect 6354 67118 6356 67170
rect 6300 67116 6356 67118
rect 5852 66834 5908 66836
rect 5852 66782 5854 66834
rect 5854 66782 5906 66834
rect 5906 66782 5908 66834
rect 5852 66780 5908 66782
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 59612 67900 59668 67956
rect 60060 67954 60116 67956
rect 60060 67902 60062 67954
rect 60062 67902 60114 67954
rect 60114 67902 60116 67954
rect 60060 67900 60116 67902
rect 81276 131738 81332 131740
rect 81276 131686 81278 131738
rect 81278 131686 81330 131738
rect 81330 131686 81332 131738
rect 81276 131684 81332 131686
rect 81380 131738 81436 131740
rect 81380 131686 81382 131738
rect 81382 131686 81434 131738
rect 81434 131686 81436 131738
rect 81380 131684 81436 131686
rect 81484 131738 81540 131740
rect 81484 131686 81486 131738
rect 81486 131686 81538 131738
rect 81538 131686 81540 131738
rect 81484 131684 81540 131686
rect 111996 131738 112052 131740
rect 111996 131686 111998 131738
rect 111998 131686 112050 131738
rect 112050 131686 112052 131738
rect 111996 131684 112052 131686
rect 112100 131738 112156 131740
rect 112100 131686 112102 131738
rect 112102 131686 112154 131738
rect 112154 131686 112156 131738
rect 112100 131684 112156 131686
rect 112204 131738 112260 131740
rect 112204 131686 112206 131738
rect 112206 131686 112258 131738
rect 112258 131686 112260 131738
rect 112204 131684 112260 131686
rect 65916 130954 65972 130956
rect 65916 130902 65918 130954
rect 65918 130902 65970 130954
rect 65970 130902 65972 130954
rect 65916 130900 65972 130902
rect 66020 130954 66076 130956
rect 66020 130902 66022 130954
rect 66022 130902 66074 130954
rect 66074 130902 66076 130954
rect 66020 130900 66076 130902
rect 66124 130954 66180 130956
rect 66124 130902 66126 130954
rect 66126 130902 66178 130954
rect 66178 130902 66180 130954
rect 66124 130900 66180 130902
rect 96636 130954 96692 130956
rect 96636 130902 96638 130954
rect 96638 130902 96690 130954
rect 96690 130902 96692 130954
rect 96636 130900 96692 130902
rect 96740 130954 96796 130956
rect 96740 130902 96742 130954
rect 96742 130902 96794 130954
rect 96794 130902 96796 130954
rect 96740 130900 96796 130902
rect 96844 130954 96900 130956
rect 96844 130902 96846 130954
rect 96846 130902 96898 130954
rect 96898 130902 96900 130954
rect 96844 130900 96900 130902
rect 81276 130170 81332 130172
rect 81276 130118 81278 130170
rect 81278 130118 81330 130170
rect 81330 130118 81332 130170
rect 81276 130116 81332 130118
rect 81380 130170 81436 130172
rect 81380 130118 81382 130170
rect 81382 130118 81434 130170
rect 81434 130118 81436 130170
rect 81380 130116 81436 130118
rect 81484 130170 81540 130172
rect 81484 130118 81486 130170
rect 81486 130118 81538 130170
rect 81538 130118 81540 130170
rect 81484 130116 81540 130118
rect 111996 130170 112052 130172
rect 111996 130118 111998 130170
rect 111998 130118 112050 130170
rect 112050 130118 112052 130170
rect 111996 130116 112052 130118
rect 112100 130170 112156 130172
rect 112100 130118 112102 130170
rect 112102 130118 112154 130170
rect 112154 130118 112156 130170
rect 112100 130116 112156 130118
rect 112204 130170 112260 130172
rect 112204 130118 112206 130170
rect 112206 130118 112258 130170
rect 112258 130118 112260 130170
rect 112204 130116 112260 130118
rect 65916 129386 65972 129388
rect 65916 129334 65918 129386
rect 65918 129334 65970 129386
rect 65970 129334 65972 129386
rect 65916 129332 65972 129334
rect 66020 129386 66076 129388
rect 66020 129334 66022 129386
rect 66022 129334 66074 129386
rect 66074 129334 66076 129386
rect 66020 129332 66076 129334
rect 66124 129386 66180 129388
rect 66124 129334 66126 129386
rect 66126 129334 66178 129386
rect 66178 129334 66180 129386
rect 66124 129332 66180 129334
rect 96636 129386 96692 129388
rect 96636 129334 96638 129386
rect 96638 129334 96690 129386
rect 96690 129334 96692 129386
rect 96636 129332 96692 129334
rect 96740 129386 96796 129388
rect 96740 129334 96742 129386
rect 96742 129334 96794 129386
rect 96794 129334 96796 129386
rect 96740 129332 96796 129334
rect 96844 129386 96900 129388
rect 96844 129334 96846 129386
rect 96846 129334 96898 129386
rect 96898 129334 96900 129386
rect 96844 129332 96900 129334
rect 81276 128602 81332 128604
rect 81276 128550 81278 128602
rect 81278 128550 81330 128602
rect 81330 128550 81332 128602
rect 81276 128548 81332 128550
rect 81380 128602 81436 128604
rect 81380 128550 81382 128602
rect 81382 128550 81434 128602
rect 81434 128550 81436 128602
rect 81380 128548 81436 128550
rect 81484 128602 81540 128604
rect 81484 128550 81486 128602
rect 81486 128550 81538 128602
rect 81538 128550 81540 128602
rect 81484 128548 81540 128550
rect 111996 128602 112052 128604
rect 111996 128550 111998 128602
rect 111998 128550 112050 128602
rect 112050 128550 112052 128602
rect 111996 128548 112052 128550
rect 112100 128602 112156 128604
rect 112100 128550 112102 128602
rect 112102 128550 112154 128602
rect 112154 128550 112156 128602
rect 112100 128548 112156 128550
rect 112204 128602 112260 128604
rect 112204 128550 112206 128602
rect 112206 128550 112258 128602
rect 112258 128550 112260 128602
rect 112204 128548 112260 128550
rect 65916 127818 65972 127820
rect 65916 127766 65918 127818
rect 65918 127766 65970 127818
rect 65970 127766 65972 127818
rect 65916 127764 65972 127766
rect 66020 127818 66076 127820
rect 66020 127766 66022 127818
rect 66022 127766 66074 127818
rect 66074 127766 66076 127818
rect 66020 127764 66076 127766
rect 66124 127818 66180 127820
rect 66124 127766 66126 127818
rect 66126 127766 66178 127818
rect 66178 127766 66180 127818
rect 66124 127764 66180 127766
rect 96636 127818 96692 127820
rect 96636 127766 96638 127818
rect 96638 127766 96690 127818
rect 96690 127766 96692 127818
rect 96636 127764 96692 127766
rect 96740 127818 96796 127820
rect 96740 127766 96742 127818
rect 96742 127766 96794 127818
rect 96794 127766 96796 127818
rect 96740 127764 96796 127766
rect 96844 127818 96900 127820
rect 96844 127766 96846 127818
rect 96846 127766 96898 127818
rect 96898 127766 96900 127818
rect 96844 127764 96900 127766
rect 81276 127034 81332 127036
rect 81276 126982 81278 127034
rect 81278 126982 81330 127034
rect 81330 126982 81332 127034
rect 81276 126980 81332 126982
rect 81380 127034 81436 127036
rect 81380 126982 81382 127034
rect 81382 126982 81434 127034
rect 81434 126982 81436 127034
rect 81380 126980 81436 126982
rect 81484 127034 81540 127036
rect 81484 126982 81486 127034
rect 81486 126982 81538 127034
rect 81538 126982 81540 127034
rect 81484 126980 81540 126982
rect 111996 127034 112052 127036
rect 111996 126982 111998 127034
rect 111998 126982 112050 127034
rect 112050 126982 112052 127034
rect 111996 126980 112052 126982
rect 112100 127034 112156 127036
rect 112100 126982 112102 127034
rect 112102 126982 112154 127034
rect 112154 126982 112156 127034
rect 112100 126980 112156 126982
rect 112204 127034 112260 127036
rect 112204 126982 112206 127034
rect 112206 126982 112258 127034
rect 112258 126982 112260 127034
rect 112204 126980 112260 126982
rect 118076 126364 118132 126420
rect 65916 126250 65972 126252
rect 65916 126198 65918 126250
rect 65918 126198 65970 126250
rect 65970 126198 65972 126250
rect 65916 126196 65972 126198
rect 66020 126250 66076 126252
rect 66020 126198 66022 126250
rect 66022 126198 66074 126250
rect 66074 126198 66076 126250
rect 66020 126196 66076 126198
rect 66124 126250 66180 126252
rect 66124 126198 66126 126250
rect 66126 126198 66178 126250
rect 66178 126198 66180 126250
rect 66124 126196 66180 126198
rect 96636 126250 96692 126252
rect 96636 126198 96638 126250
rect 96638 126198 96690 126250
rect 96690 126198 96692 126250
rect 96636 126196 96692 126198
rect 96740 126250 96796 126252
rect 96740 126198 96742 126250
rect 96742 126198 96794 126250
rect 96794 126198 96796 126250
rect 96740 126196 96796 126198
rect 96844 126250 96900 126252
rect 96844 126198 96846 126250
rect 96846 126198 96898 126250
rect 96898 126198 96900 126250
rect 96844 126196 96900 126198
rect 81276 125466 81332 125468
rect 81276 125414 81278 125466
rect 81278 125414 81330 125466
rect 81330 125414 81332 125466
rect 81276 125412 81332 125414
rect 81380 125466 81436 125468
rect 81380 125414 81382 125466
rect 81382 125414 81434 125466
rect 81434 125414 81436 125466
rect 81380 125412 81436 125414
rect 81484 125466 81540 125468
rect 81484 125414 81486 125466
rect 81486 125414 81538 125466
rect 81538 125414 81540 125466
rect 81484 125412 81540 125414
rect 111996 125466 112052 125468
rect 111996 125414 111998 125466
rect 111998 125414 112050 125466
rect 112050 125414 112052 125466
rect 111996 125412 112052 125414
rect 112100 125466 112156 125468
rect 112100 125414 112102 125466
rect 112102 125414 112154 125466
rect 112154 125414 112156 125466
rect 112100 125412 112156 125414
rect 112204 125466 112260 125468
rect 112204 125414 112206 125466
rect 112206 125414 112258 125466
rect 112258 125414 112260 125466
rect 112204 125412 112260 125414
rect 65916 124682 65972 124684
rect 65916 124630 65918 124682
rect 65918 124630 65970 124682
rect 65970 124630 65972 124682
rect 65916 124628 65972 124630
rect 66020 124682 66076 124684
rect 66020 124630 66022 124682
rect 66022 124630 66074 124682
rect 66074 124630 66076 124682
rect 66020 124628 66076 124630
rect 66124 124682 66180 124684
rect 66124 124630 66126 124682
rect 66126 124630 66178 124682
rect 66178 124630 66180 124682
rect 66124 124628 66180 124630
rect 96636 124682 96692 124684
rect 96636 124630 96638 124682
rect 96638 124630 96690 124682
rect 96690 124630 96692 124682
rect 96636 124628 96692 124630
rect 96740 124682 96796 124684
rect 96740 124630 96742 124682
rect 96742 124630 96794 124682
rect 96794 124630 96796 124682
rect 96740 124628 96796 124630
rect 96844 124682 96900 124684
rect 96844 124630 96846 124682
rect 96846 124630 96898 124682
rect 96898 124630 96900 124682
rect 96844 124628 96900 124630
rect 81276 123898 81332 123900
rect 81276 123846 81278 123898
rect 81278 123846 81330 123898
rect 81330 123846 81332 123898
rect 81276 123844 81332 123846
rect 81380 123898 81436 123900
rect 81380 123846 81382 123898
rect 81382 123846 81434 123898
rect 81434 123846 81436 123898
rect 81380 123844 81436 123846
rect 81484 123898 81540 123900
rect 81484 123846 81486 123898
rect 81486 123846 81538 123898
rect 81538 123846 81540 123898
rect 81484 123844 81540 123846
rect 111996 123898 112052 123900
rect 111996 123846 111998 123898
rect 111998 123846 112050 123898
rect 112050 123846 112052 123898
rect 111996 123844 112052 123846
rect 112100 123898 112156 123900
rect 112100 123846 112102 123898
rect 112102 123846 112154 123898
rect 112154 123846 112156 123898
rect 112100 123844 112156 123846
rect 112204 123898 112260 123900
rect 112204 123846 112206 123898
rect 112206 123846 112258 123898
rect 112258 123846 112260 123898
rect 112204 123844 112260 123846
rect 118076 123676 118132 123732
rect 65916 123114 65972 123116
rect 65916 123062 65918 123114
rect 65918 123062 65970 123114
rect 65970 123062 65972 123114
rect 65916 123060 65972 123062
rect 66020 123114 66076 123116
rect 66020 123062 66022 123114
rect 66022 123062 66074 123114
rect 66074 123062 66076 123114
rect 66020 123060 66076 123062
rect 66124 123114 66180 123116
rect 66124 123062 66126 123114
rect 66126 123062 66178 123114
rect 66178 123062 66180 123114
rect 66124 123060 66180 123062
rect 96636 123114 96692 123116
rect 96636 123062 96638 123114
rect 96638 123062 96690 123114
rect 96690 123062 96692 123114
rect 96636 123060 96692 123062
rect 96740 123114 96796 123116
rect 96740 123062 96742 123114
rect 96742 123062 96794 123114
rect 96794 123062 96796 123114
rect 96740 123060 96796 123062
rect 96844 123114 96900 123116
rect 96844 123062 96846 123114
rect 96846 123062 96898 123114
rect 96898 123062 96900 123114
rect 96844 123060 96900 123062
rect 81276 122330 81332 122332
rect 81276 122278 81278 122330
rect 81278 122278 81330 122330
rect 81330 122278 81332 122330
rect 81276 122276 81332 122278
rect 81380 122330 81436 122332
rect 81380 122278 81382 122330
rect 81382 122278 81434 122330
rect 81434 122278 81436 122330
rect 81380 122276 81436 122278
rect 81484 122330 81540 122332
rect 81484 122278 81486 122330
rect 81486 122278 81538 122330
rect 81538 122278 81540 122330
rect 81484 122276 81540 122278
rect 111996 122330 112052 122332
rect 111996 122278 111998 122330
rect 111998 122278 112050 122330
rect 112050 122278 112052 122330
rect 111996 122276 112052 122278
rect 112100 122330 112156 122332
rect 112100 122278 112102 122330
rect 112102 122278 112154 122330
rect 112154 122278 112156 122330
rect 112100 122276 112156 122278
rect 112204 122330 112260 122332
rect 112204 122278 112206 122330
rect 112206 122278 112258 122330
rect 112258 122278 112260 122330
rect 112204 122276 112260 122278
rect 65916 121546 65972 121548
rect 65916 121494 65918 121546
rect 65918 121494 65970 121546
rect 65970 121494 65972 121546
rect 65916 121492 65972 121494
rect 66020 121546 66076 121548
rect 66020 121494 66022 121546
rect 66022 121494 66074 121546
rect 66074 121494 66076 121546
rect 66020 121492 66076 121494
rect 66124 121546 66180 121548
rect 66124 121494 66126 121546
rect 66126 121494 66178 121546
rect 66178 121494 66180 121546
rect 66124 121492 66180 121494
rect 96636 121546 96692 121548
rect 96636 121494 96638 121546
rect 96638 121494 96690 121546
rect 96690 121494 96692 121546
rect 96636 121492 96692 121494
rect 96740 121546 96796 121548
rect 96740 121494 96742 121546
rect 96742 121494 96794 121546
rect 96794 121494 96796 121546
rect 96740 121492 96796 121494
rect 96844 121546 96900 121548
rect 96844 121494 96846 121546
rect 96846 121494 96898 121546
rect 96898 121494 96900 121546
rect 96844 121492 96900 121494
rect 81276 120762 81332 120764
rect 81276 120710 81278 120762
rect 81278 120710 81330 120762
rect 81330 120710 81332 120762
rect 81276 120708 81332 120710
rect 81380 120762 81436 120764
rect 81380 120710 81382 120762
rect 81382 120710 81434 120762
rect 81434 120710 81436 120762
rect 81380 120708 81436 120710
rect 81484 120762 81540 120764
rect 81484 120710 81486 120762
rect 81486 120710 81538 120762
rect 81538 120710 81540 120762
rect 81484 120708 81540 120710
rect 111996 120762 112052 120764
rect 111996 120710 111998 120762
rect 111998 120710 112050 120762
rect 112050 120710 112052 120762
rect 111996 120708 112052 120710
rect 112100 120762 112156 120764
rect 112100 120710 112102 120762
rect 112102 120710 112154 120762
rect 112154 120710 112156 120762
rect 112100 120708 112156 120710
rect 112204 120762 112260 120764
rect 112204 120710 112206 120762
rect 112206 120710 112258 120762
rect 112258 120710 112260 120762
rect 112204 120708 112260 120710
rect 65916 119978 65972 119980
rect 65916 119926 65918 119978
rect 65918 119926 65970 119978
rect 65970 119926 65972 119978
rect 65916 119924 65972 119926
rect 66020 119978 66076 119980
rect 66020 119926 66022 119978
rect 66022 119926 66074 119978
rect 66074 119926 66076 119978
rect 66020 119924 66076 119926
rect 66124 119978 66180 119980
rect 66124 119926 66126 119978
rect 66126 119926 66178 119978
rect 66178 119926 66180 119978
rect 66124 119924 66180 119926
rect 96636 119978 96692 119980
rect 96636 119926 96638 119978
rect 96638 119926 96690 119978
rect 96690 119926 96692 119978
rect 96636 119924 96692 119926
rect 96740 119978 96796 119980
rect 96740 119926 96742 119978
rect 96742 119926 96794 119978
rect 96794 119926 96796 119978
rect 96740 119924 96796 119926
rect 96844 119978 96900 119980
rect 96844 119926 96846 119978
rect 96846 119926 96898 119978
rect 96898 119926 96900 119978
rect 96844 119924 96900 119926
rect 81276 119194 81332 119196
rect 81276 119142 81278 119194
rect 81278 119142 81330 119194
rect 81330 119142 81332 119194
rect 81276 119140 81332 119142
rect 81380 119194 81436 119196
rect 81380 119142 81382 119194
rect 81382 119142 81434 119194
rect 81434 119142 81436 119194
rect 81380 119140 81436 119142
rect 81484 119194 81540 119196
rect 81484 119142 81486 119194
rect 81486 119142 81538 119194
rect 81538 119142 81540 119194
rect 81484 119140 81540 119142
rect 111996 119194 112052 119196
rect 111996 119142 111998 119194
rect 111998 119142 112050 119194
rect 112050 119142 112052 119194
rect 111996 119140 112052 119142
rect 112100 119194 112156 119196
rect 112100 119142 112102 119194
rect 112102 119142 112154 119194
rect 112154 119142 112156 119194
rect 112100 119140 112156 119142
rect 112204 119194 112260 119196
rect 112204 119142 112206 119194
rect 112206 119142 112258 119194
rect 112258 119142 112260 119194
rect 112204 119140 112260 119142
rect 65916 118410 65972 118412
rect 65916 118358 65918 118410
rect 65918 118358 65970 118410
rect 65970 118358 65972 118410
rect 65916 118356 65972 118358
rect 66020 118410 66076 118412
rect 66020 118358 66022 118410
rect 66022 118358 66074 118410
rect 66074 118358 66076 118410
rect 66020 118356 66076 118358
rect 66124 118410 66180 118412
rect 66124 118358 66126 118410
rect 66126 118358 66178 118410
rect 66178 118358 66180 118410
rect 66124 118356 66180 118358
rect 96636 118410 96692 118412
rect 96636 118358 96638 118410
rect 96638 118358 96690 118410
rect 96690 118358 96692 118410
rect 96636 118356 96692 118358
rect 96740 118410 96796 118412
rect 96740 118358 96742 118410
rect 96742 118358 96794 118410
rect 96794 118358 96796 118410
rect 96740 118356 96796 118358
rect 96844 118410 96900 118412
rect 96844 118358 96846 118410
rect 96846 118358 96898 118410
rect 96898 118358 96900 118410
rect 96844 118356 96900 118358
rect 81276 117626 81332 117628
rect 81276 117574 81278 117626
rect 81278 117574 81330 117626
rect 81330 117574 81332 117626
rect 81276 117572 81332 117574
rect 81380 117626 81436 117628
rect 81380 117574 81382 117626
rect 81382 117574 81434 117626
rect 81434 117574 81436 117626
rect 81380 117572 81436 117574
rect 81484 117626 81540 117628
rect 81484 117574 81486 117626
rect 81486 117574 81538 117626
rect 81538 117574 81540 117626
rect 81484 117572 81540 117574
rect 111996 117626 112052 117628
rect 111996 117574 111998 117626
rect 111998 117574 112050 117626
rect 112050 117574 112052 117626
rect 111996 117572 112052 117574
rect 112100 117626 112156 117628
rect 112100 117574 112102 117626
rect 112102 117574 112154 117626
rect 112154 117574 112156 117626
rect 112100 117572 112156 117574
rect 112204 117626 112260 117628
rect 112204 117574 112206 117626
rect 112206 117574 112258 117626
rect 112258 117574 112260 117626
rect 112204 117572 112260 117574
rect 65916 116842 65972 116844
rect 65916 116790 65918 116842
rect 65918 116790 65970 116842
rect 65970 116790 65972 116842
rect 65916 116788 65972 116790
rect 66020 116842 66076 116844
rect 66020 116790 66022 116842
rect 66022 116790 66074 116842
rect 66074 116790 66076 116842
rect 66020 116788 66076 116790
rect 66124 116842 66180 116844
rect 66124 116790 66126 116842
rect 66126 116790 66178 116842
rect 66178 116790 66180 116842
rect 66124 116788 66180 116790
rect 96636 116842 96692 116844
rect 96636 116790 96638 116842
rect 96638 116790 96690 116842
rect 96690 116790 96692 116842
rect 96636 116788 96692 116790
rect 96740 116842 96796 116844
rect 96740 116790 96742 116842
rect 96742 116790 96794 116842
rect 96794 116790 96796 116842
rect 96740 116788 96796 116790
rect 96844 116842 96900 116844
rect 96844 116790 96846 116842
rect 96846 116790 96898 116842
rect 96898 116790 96900 116842
rect 96844 116788 96900 116790
rect 118076 116338 118132 116340
rect 118076 116286 118078 116338
rect 118078 116286 118130 116338
rect 118130 116286 118132 116338
rect 118076 116284 118132 116286
rect 81276 116058 81332 116060
rect 81276 116006 81278 116058
rect 81278 116006 81330 116058
rect 81330 116006 81332 116058
rect 81276 116004 81332 116006
rect 81380 116058 81436 116060
rect 81380 116006 81382 116058
rect 81382 116006 81434 116058
rect 81434 116006 81436 116058
rect 81380 116004 81436 116006
rect 81484 116058 81540 116060
rect 81484 116006 81486 116058
rect 81486 116006 81538 116058
rect 81538 116006 81540 116058
rect 81484 116004 81540 116006
rect 111996 116058 112052 116060
rect 111996 116006 111998 116058
rect 111998 116006 112050 116058
rect 112050 116006 112052 116058
rect 111996 116004 112052 116006
rect 112100 116058 112156 116060
rect 112100 116006 112102 116058
rect 112102 116006 112154 116058
rect 112154 116006 112156 116058
rect 112100 116004 112156 116006
rect 112204 116058 112260 116060
rect 112204 116006 112206 116058
rect 112206 116006 112258 116058
rect 112258 116006 112260 116058
rect 112204 116004 112260 116006
rect 65916 115274 65972 115276
rect 65916 115222 65918 115274
rect 65918 115222 65970 115274
rect 65970 115222 65972 115274
rect 65916 115220 65972 115222
rect 66020 115274 66076 115276
rect 66020 115222 66022 115274
rect 66022 115222 66074 115274
rect 66074 115222 66076 115274
rect 66020 115220 66076 115222
rect 66124 115274 66180 115276
rect 66124 115222 66126 115274
rect 66126 115222 66178 115274
rect 66178 115222 66180 115274
rect 66124 115220 66180 115222
rect 96636 115274 96692 115276
rect 96636 115222 96638 115274
rect 96638 115222 96690 115274
rect 96690 115222 96692 115274
rect 96636 115220 96692 115222
rect 96740 115274 96796 115276
rect 96740 115222 96742 115274
rect 96742 115222 96794 115274
rect 96794 115222 96796 115274
rect 96740 115220 96796 115222
rect 96844 115274 96900 115276
rect 96844 115222 96846 115274
rect 96846 115222 96898 115274
rect 96898 115222 96900 115274
rect 96844 115220 96900 115222
rect 118076 114940 118132 114996
rect 81276 114490 81332 114492
rect 81276 114438 81278 114490
rect 81278 114438 81330 114490
rect 81330 114438 81332 114490
rect 81276 114436 81332 114438
rect 81380 114490 81436 114492
rect 81380 114438 81382 114490
rect 81382 114438 81434 114490
rect 81434 114438 81436 114490
rect 81380 114436 81436 114438
rect 81484 114490 81540 114492
rect 81484 114438 81486 114490
rect 81486 114438 81538 114490
rect 81538 114438 81540 114490
rect 81484 114436 81540 114438
rect 111996 114490 112052 114492
rect 111996 114438 111998 114490
rect 111998 114438 112050 114490
rect 112050 114438 112052 114490
rect 111996 114436 112052 114438
rect 112100 114490 112156 114492
rect 112100 114438 112102 114490
rect 112102 114438 112154 114490
rect 112154 114438 112156 114490
rect 112100 114436 112156 114438
rect 112204 114490 112260 114492
rect 112204 114438 112206 114490
rect 112206 114438 112258 114490
rect 112258 114438 112260 114490
rect 112204 114436 112260 114438
rect 65916 113706 65972 113708
rect 65916 113654 65918 113706
rect 65918 113654 65970 113706
rect 65970 113654 65972 113706
rect 65916 113652 65972 113654
rect 66020 113706 66076 113708
rect 66020 113654 66022 113706
rect 66022 113654 66074 113706
rect 66074 113654 66076 113706
rect 66020 113652 66076 113654
rect 66124 113706 66180 113708
rect 66124 113654 66126 113706
rect 66126 113654 66178 113706
rect 66178 113654 66180 113706
rect 66124 113652 66180 113654
rect 96636 113706 96692 113708
rect 96636 113654 96638 113706
rect 96638 113654 96690 113706
rect 96690 113654 96692 113706
rect 96636 113652 96692 113654
rect 96740 113706 96796 113708
rect 96740 113654 96742 113706
rect 96742 113654 96794 113706
rect 96794 113654 96796 113706
rect 96740 113652 96796 113654
rect 96844 113706 96900 113708
rect 96844 113654 96846 113706
rect 96846 113654 96898 113706
rect 96898 113654 96900 113706
rect 96844 113652 96900 113654
rect 117628 113596 117684 113652
rect 81276 112922 81332 112924
rect 81276 112870 81278 112922
rect 81278 112870 81330 112922
rect 81330 112870 81332 112922
rect 81276 112868 81332 112870
rect 81380 112922 81436 112924
rect 81380 112870 81382 112922
rect 81382 112870 81434 112922
rect 81434 112870 81436 112922
rect 81380 112868 81436 112870
rect 81484 112922 81540 112924
rect 81484 112870 81486 112922
rect 81486 112870 81538 112922
rect 81538 112870 81540 112922
rect 81484 112868 81540 112870
rect 111996 112922 112052 112924
rect 111996 112870 111998 112922
rect 111998 112870 112050 112922
rect 112050 112870 112052 112922
rect 111996 112868 112052 112870
rect 112100 112922 112156 112924
rect 112100 112870 112102 112922
rect 112102 112870 112154 112922
rect 112154 112870 112156 112922
rect 112100 112868 112156 112870
rect 112204 112922 112260 112924
rect 112204 112870 112206 112922
rect 112206 112870 112258 112922
rect 112258 112870 112260 112922
rect 112204 112868 112260 112870
rect 65916 112138 65972 112140
rect 65916 112086 65918 112138
rect 65918 112086 65970 112138
rect 65970 112086 65972 112138
rect 65916 112084 65972 112086
rect 66020 112138 66076 112140
rect 66020 112086 66022 112138
rect 66022 112086 66074 112138
rect 66074 112086 66076 112138
rect 66020 112084 66076 112086
rect 66124 112138 66180 112140
rect 66124 112086 66126 112138
rect 66126 112086 66178 112138
rect 66178 112086 66180 112138
rect 66124 112084 66180 112086
rect 96636 112138 96692 112140
rect 96636 112086 96638 112138
rect 96638 112086 96690 112138
rect 96690 112086 96692 112138
rect 96636 112084 96692 112086
rect 96740 112138 96796 112140
rect 96740 112086 96742 112138
rect 96742 112086 96794 112138
rect 96794 112086 96796 112138
rect 96740 112084 96796 112086
rect 96844 112138 96900 112140
rect 96844 112086 96846 112138
rect 96846 112086 96898 112138
rect 96898 112086 96900 112138
rect 96844 112084 96900 112086
rect 118076 111634 118132 111636
rect 118076 111582 118078 111634
rect 118078 111582 118130 111634
rect 118130 111582 118132 111634
rect 118076 111580 118132 111582
rect 81276 111354 81332 111356
rect 81276 111302 81278 111354
rect 81278 111302 81330 111354
rect 81330 111302 81332 111354
rect 81276 111300 81332 111302
rect 81380 111354 81436 111356
rect 81380 111302 81382 111354
rect 81382 111302 81434 111354
rect 81434 111302 81436 111354
rect 81380 111300 81436 111302
rect 81484 111354 81540 111356
rect 81484 111302 81486 111354
rect 81486 111302 81538 111354
rect 81538 111302 81540 111354
rect 81484 111300 81540 111302
rect 111996 111354 112052 111356
rect 111996 111302 111998 111354
rect 111998 111302 112050 111354
rect 112050 111302 112052 111354
rect 111996 111300 112052 111302
rect 112100 111354 112156 111356
rect 112100 111302 112102 111354
rect 112102 111302 112154 111354
rect 112154 111302 112156 111354
rect 112100 111300 112156 111302
rect 112204 111354 112260 111356
rect 112204 111302 112206 111354
rect 112206 111302 112258 111354
rect 112258 111302 112260 111354
rect 112204 111300 112260 111302
rect 65916 110570 65972 110572
rect 65916 110518 65918 110570
rect 65918 110518 65970 110570
rect 65970 110518 65972 110570
rect 65916 110516 65972 110518
rect 66020 110570 66076 110572
rect 66020 110518 66022 110570
rect 66022 110518 66074 110570
rect 66074 110518 66076 110570
rect 66020 110516 66076 110518
rect 66124 110570 66180 110572
rect 66124 110518 66126 110570
rect 66126 110518 66178 110570
rect 66178 110518 66180 110570
rect 66124 110516 66180 110518
rect 96636 110570 96692 110572
rect 96636 110518 96638 110570
rect 96638 110518 96690 110570
rect 96690 110518 96692 110570
rect 96636 110516 96692 110518
rect 96740 110570 96796 110572
rect 96740 110518 96742 110570
rect 96742 110518 96794 110570
rect 96794 110518 96796 110570
rect 96740 110516 96796 110518
rect 96844 110570 96900 110572
rect 96844 110518 96846 110570
rect 96846 110518 96898 110570
rect 96898 110518 96900 110570
rect 96844 110516 96900 110518
rect 118076 110236 118132 110292
rect 81276 109786 81332 109788
rect 81276 109734 81278 109786
rect 81278 109734 81330 109786
rect 81330 109734 81332 109786
rect 81276 109732 81332 109734
rect 81380 109786 81436 109788
rect 81380 109734 81382 109786
rect 81382 109734 81434 109786
rect 81434 109734 81436 109786
rect 81380 109732 81436 109734
rect 81484 109786 81540 109788
rect 81484 109734 81486 109786
rect 81486 109734 81538 109786
rect 81538 109734 81540 109786
rect 81484 109732 81540 109734
rect 111996 109786 112052 109788
rect 111996 109734 111998 109786
rect 111998 109734 112050 109786
rect 112050 109734 112052 109786
rect 111996 109732 112052 109734
rect 112100 109786 112156 109788
rect 112100 109734 112102 109786
rect 112102 109734 112154 109786
rect 112154 109734 112156 109786
rect 112100 109732 112156 109734
rect 112204 109786 112260 109788
rect 112204 109734 112206 109786
rect 112206 109734 112258 109786
rect 112258 109734 112260 109786
rect 112204 109732 112260 109734
rect 65916 109002 65972 109004
rect 65916 108950 65918 109002
rect 65918 108950 65970 109002
rect 65970 108950 65972 109002
rect 65916 108948 65972 108950
rect 66020 109002 66076 109004
rect 66020 108950 66022 109002
rect 66022 108950 66074 109002
rect 66074 108950 66076 109002
rect 66020 108948 66076 108950
rect 66124 109002 66180 109004
rect 66124 108950 66126 109002
rect 66126 108950 66178 109002
rect 66178 108950 66180 109002
rect 66124 108948 66180 108950
rect 96636 109002 96692 109004
rect 96636 108950 96638 109002
rect 96638 108950 96690 109002
rect 96690 108950 96692 109002
rect 96636 108948 96692 108950
rect 96740 109002 96796 109004
rect 96740 108950 96742 109002
rect 96742 108950 96794 109002
rect 96794 108950 96796 109002
rect 96740 108948 96796 108950
rect 96844 109002 96900 109004
rect 96844 108950 96846 109002
rect 96846 108950 96898 109002
rect 96898 108950 96900 109002
rect 96844 108948 96900 108950
rect 81276 108218 81332 108220
rect 81276 108166 81278 108218
rect 81278 108166 81330 108218
rect 81330 108166 81332 108218
rect 81276 108164 81332 108166
rect 81380 108218 81436 108220
rect 81380 108166 81382 108218
rect 81382 108166 81434 108218
rect 81434 108166 81436 108218
rect 81380 108164 81436 108166
rect 81484 108218 81540 108220
rect 81484 108166 81486 108218
rect 81486 108166 81538 108218
rect 81538 108166 81540 108218
rect 81484 108164 81540 108166
rect 111996 108218 112052 108220
rect 111996 108166 111998 108218
rect 111998 108166 112050 108218
rect 112050 108166 112052 108218
rect 111996 108164 112052 108166
rect 112100 108218 112156 108220
rect 112100 108166 112102 108218
rect 112102 108166 112154 108218
rect 112154 108166 112156 108218
rect 112100 108164 112156 108166
rect 112204 108218 112260 108220
rect 112204 108166 112206 108218
rect 112206 108166 112258 108218
rect 112258 108166 112260 108218
rect 112204 108164 112260 108166
rect 118076 107548 118132 107604
rect 65916 107434 65972 107436
rect 65916 107382 65918 107434
rect 65918 107382 65970 107434
rect 65970 107382 65972 107434
rect 65916 107380 65972 107382
rect 66020 107434 66076 107436
rect 66020 107382 66022 107434
rect 66022 107382 66074 107434
rect 66074 107382 66076 107434
rect 66020 107380 66076 107382
rect 66124 107434 66180 107436
rect 66124 107382 66126 107434
rect 66126 107382 66178 107434
rect 66178 107382 66180 107434
rect 66124 107380 66180 107382
rect 96636 107434 96692 107436
rect 96636 107382 96638 107434
rect 96638 107382 96690 107434
rect 96690 107382 96692 107434
rect 96636 107380 96692 107382
rect 96740 107434 96796 107436
rect 96740 107382 96742 107434
rect 96742 107382 96794 107434
rect 96794 107382 96796 107434
rect 96740 107380 96796 107382
rect 96844 107434 96900 107436
rect 96844 107382 96846 107434
rect 96846 107382 96898 107434
rect 96898 107382 96900 107434
rect 96844 107380 96900 107382
rect 81276 106650 81332 106652
rect 81276 106598 81278 106650
rect 81278 106598 81330 106650
rect 81330 106598 81332 106650
rect 81276 106596 81332 106598
rect 81380 106650 81436 106652
rect 81380 106598 81382 106650
rect 81382 106598 81434 106650
rect 81434 106598 81436 106650
rect 81380 106596 81436 106598
rect 81484 106650 81540 106652
rect 81484 106598 81486 106650
rect 81486 106598 81538 106650
rect 81538 106598 81540 106650
rect 81484 106596 81540 106598
rect 111996 106650 112052 106652
rect 111996 106598 111998 106650
rect 111998 106598 112050 106650
rect 112050 106598 112052 106650
rect 111996 106596 112052 106598
rect 112100 106650 112156 106652
rect 112100 106598 112102 106650
rect 112102 106598 112154 106650
rect 112154 106598 112156 106650
rect 112100 106596 112156 106598
rect 112204 106650 112260 106652
rect 112204 106598 112206 106650
rect 112206 106598 112258 106650
rect 112258 106598 112260 106650
rect 112204 106596 112260 106598
rect 118076 106204 118132 106260
rect 65916 105866 65972 105868
rect 65916 105814 65918 105866
rect 65918 105814 65970 105866
rect 65970 105814 65972 105866
rect 65916 105812 65972 105814
rect 66020 105866 66076 105868
rect 66020 105814 66022 105866
rect 66022 105814 66074 105866
rect 66074 105814 66076 105866
rect 66020 105812 66076 105814
rect 66124 105866 66180 105868
rect 66124 105814 66126 105866
rect 66126 105814 66178 105866
rect 66178 105814 66180 105866
rect 66124 105812 66180 105814
rect 96636 105866 96692 105868
rect 96636 105814 96638 105866
rect 96638 105814 96690 105866
rect 96690 105814 96692 105866
rect 96636 105812 96692 105814
rect 96740 105866 96796 105868
rect 96740 105814 96742 105866
rect 96742 105814 96794 105866
rect 96794 105814 96796 105866
rect 96740 105812 96796 105814
rect 96844 105866 96900 105868
rect 96844 105814 96846 105866
rect 96846 105814 96898 105866
rect 96898 105814 96900 105866
rect 96844 105812 96900 105814
rect 81276 105082 81332 105084
rect 81276 105030 81278 105082
rect 81278 105030 81330 105082
rect 81330 105030 81332 105082
rect 81276 105028 81332 105030
rect 81380 105082 81436 105084
rect 81380 105030 81382 105082
rect 81382 105030 81434 105082
rect 81434 105030 81436 105082
rect 81380 105028 81436 105030
rect 81484 105082 81540 105084
rect 81484 105030 81486 105082
rect 81486 105030 81538 105082
rect 81538 105030 81540 105082
rect 81484 105028 81540 105030
rect 111996 105082 112052 105084
rect 111996 105030 111998 105082
rect 111998 105030 112050 105082
rect 112050 105030 112052 105082
rect 111996 105028 112052 105030
rect 112100 105082 112156 105084
rect 112100 105030 112102 105082
rect 112102 105030 112154 105082
rect 112154 105030 112156 105082
rect 112100 105028 112156 105030
rect 112204 105082 112260 105084
rect 112204 105030 112206 105082
rect 112206 105030 112258 105082
rect 112258 105030 112260 105082
rect 112204 105028 112260 105030
rect 65916 104298 65972 104300
rect 65916 104246 65918 104298
rect 65918 104246 65970 104298
rect 65970 104246 65972 104298
rect 65916 104244 65972 104246
rect 66020 104298 66076 104300
rect 66020 104246 66022 104298
rect 66022 104246 66074 104298
rect 66074 104246 66076 104298
rect 66020 104244 66076 104246
rect 66124 104298 66180 104300
rect 66124 104246 66126 104298
rect 66126 104246 66178 104298
rect 66178 104246 66180 104298
rect 66124 104244 66180 104246
rect 96636 104298 96692 104300
rect 96636 104246 96638 104298
rect 96638 104246 96690 104298
rect 96690 104246 96692 104298
rect 96636 104244 96692 104246
rect 96740 104298 96796 104300
rect 96740 104246 96742 104298
rect 96742 104246 96794 104298
rect 96794 104246 96796 104298
rect 96740 104244 96796 104246
rect 96844 104298 96900 104300
rect 96844 104246 96846 104298
rect 96846 104246 96898 104298
rect 96898 104246 96900 104298
rect 96844 104244 96900 104246
rect 81276 103514 81332 103516
rect 81276 103462 81278 103514
rect 81278 103462 81330 103514
rect 81330 103462 81332 103514
rect 81276 103460 81332 103462
rect 81380 103514 81436 103516
rect 81380 103462 81382 103514
rect 81382 103462 81434 103514
rect 81434 103462 81436 103514
rect 81380 103460 81436 103462
rect 81484 103514 81540 103516
rect 81484 103462 81486 103514
rect 81486 103462 81538 103514
rect 81538 103462 81540 103514
rect 81484 103460 81540 103462
rect 111996 103514 112052 103516
rect 111996 103462 111998 103514
rect 111998 103462 112050 103514
rect 112050 103462 112052 103514
rect 111996 103460 112052 103462
rect 112100 103514 112156 103516
rect 112100 103462 112102 103514
rect 112102 103462 112154 103514
rect 112154 103462 112156 103514
rect 112100 103460 112156 103462
rect 112204 103514 112260 103516
rect 112204 103462 112206 103514
rect 112206 103462 112258 103514
rect 112258 103462 112260 103514
rect 112204 103460 112260 103462
rect 118076 102844 118132 102900
rect 65916 102730 65972 102732
rect 65916 102678 65918 102730
rect 65918 102678 65970 102730
rect 65970 102678 65972 102730
rect 65916 102676 65972 102678
rect 66020 102730 66076 102732
rect 66020 102678 66022 102730
rect 66022 102678 66074 102730
rect 66074 102678 66076 102730
rect 66020 102676 66076 102678
rect 66124 102730 66180 102732
rect 66124 102678 66126 102730
rect 66126 102678 66178 102730
rect 66178 102678 66180 102730
rect 66124 102676 66180 102678
rect 96636 102730 96692 102732
rect 96636 102678 96638 102730
rect 96638 102678 96690 102730
rect 96690 102678 96692 102730
rect 96636 102676 96692 102678
rect 96740 102730 96796 102732
rect 96740 102678 96742 102730
rect 96742 102678 96794 102730
rect 96794 102678 96796 102730
rect 96740 102676 96796 102678
rect 96844 102730 96900 102732
rect 96844 102678 96846 102730
rect 96846 102678 96898 102730
rect 96898 102678 96900 102730
rect 96844 102676 96900 102678
rect 81276 101946 81332 101948
rect 81276 101894 81278 101946
rect 81278 101894 81330 101946
rect 81330 101894 81332 101946
rect 81276 101892 81332 101894
rect 81380 101946 81436 101948
rect 81380 101894 81382 101946
rect 81382 101894 81434 101946
rect 81434 101894 81436 101946
rect 81380 101892 81436 101894
rect 81484 101946 81540 101948
rect 81484 101894 81486 101946
rect 81486 101894 81538 101946
rect 81538 101894 81540 101946
rect 81484 101892 81540 101894
rect 111996 101946 112052 101948
rect 111996 101894 111998 101946
rect 111998 101894 112050 101946
rect 112050 101894 112052 101946
rect 111996 101892 112052 101894
rect 112100 101946 112156 101948
rect 112100 101894 112102 101946
rect 112102 101894 112154 101946
rect 112154 101894 112156 101946
rect 112100 101892 112156 101894
rect 112204 101946 112260 101948
rect 112204 101894 112206 101946
rect 112206 101894 112258 101946
rect 112258 101894 112260 101946
rect 112204 101892 112260 101894
rect 65916 101162 65972 101164
rect 65916 101110 65918 101162
rect 65918 101110 65970 101162
rect 65970 101110 65972 101162
rect 65916 101108 65972 101110
rect 66020 101162 66076 101164
rect 66020 101110 66022 101162
rect 66022 101110 66074 101162
rect 66074 101110 66076 101162
rect 66020 101108 66076 101110
rect 66124 101162 66180 101164
rect 66124 101110 66126 101162
rect 66126 101110 66178 101162
rect 66178 101110 66180 101162
rect 66124 101108 66180 101110
rect 96636 101162 96692 101164
rect 96636 101110 96638 101162
rect 96638 101110 96690 101162
rect 96690 101110 96692 101162
rect 96636 101108 96692 101110
rect 96740 101162 96796 101164
rect 96740 101110 96742 101162
rect 96742 101110 96794 101162
rect 96794 101110 96796 101162
rect 96740 101108 96796 101110
rect 96844 101162 96900 101164
rect 96844 101110 96846 101162
rect 96846 101110 96898 101162
rect 96898 101110 96900 101162
rect 96844 101108 96900 101110
rect 81276 100378 81332 100380
rect 81276 100326 81278 100378
rect 81278 100326 81330 100378
rect 81330 100326 81332 100378
rect 81276 100324 81332 100326
rect 81380 100378 81436 100380
rect 81380 100326 81382 100378
rect 81382 100326 81434 100378
rect 81434 100326 81436 100378
rect 81380 100324 81436 100326
rect 81484 100378 81540 100380
rect 81484 100326 81486 100378
rect 81486 100326 81538 100378
rect 81538 100326 81540 100378
rect 81484 100324 81540 100326
rect 111996 100378 112052 100380
rect 111996 100326 111998 100378
rect 111998 100326 112050 100378
rect 112050 100326 112052 100378
rect 111996 100324 112052 100326
rect 112100 100378 112156 100380
rect 112100 100326 112102 100378
rect 112102 100326 112154 100378
rect 112154 100326 112156 100378
rect 112100 100324 112156 100326
rect 112204 100378 112260 100380
rect 112204 100326 112206 100378
rect 112206 100326 112258 100378
rect 112258 100326 112260 100378
rect 112204 100324 112260 100326
rect 65916 99594 65972 99596
rect 65916 99542 65918 99594
rect 65918 99542 65970 99594
rect 65970 99542 65972 99594
rect 65916 99540 65972 99542
rect 66020 99594 66076 99596
rect 66020 99542 66022 99594
rect 66022 99542 66074 99594
rect 66074 99542 66076 99594
rect 66020 99540 66076 99542
rect 66124 99594 66180 99596
rect 66124 99542 66126 99594
rect 66126 99542 66178 99594
rect 66178 99542 66180 99594
rect 66124 99540 66180 99542
rect 96636 99594 96692 99596
rect 96636 99542 96638 99594
rect 96638 99542 96690 99594
rect 96690 99542 96692 99594
rect 96636 99540 96692 99542
rect 96740 99594 96796 99596
rect 96740 99542 96742 99594
rect 96742 99542 96794 99594
rect 96794 99542 96796 99594
rect 96740 99540 96796 99542
rect 96844 99594 96900 99596
rect 96844 99542 96846 99594
rect 96846 99542 96898 99594
rect 96898 99542 96900 99594
rect 96844 99540 96900 99542
rect 81276 98810 81332 98812
rect 81276 98758 81278 98810
rect 81278 98758 81330 98810
rect 81330 98758 81332 98810
rect 81276 98756 81332 98758
rect 81380 98810 81436 98812
rect 81380 98758 81382 98810
rect 81382 98758 81434 98810
rect 81434 98758 81436 98810
rect 81380 98756 81436 98758
rect 81484 98810 81540 98812
rect 81484 98758 81486 98810
rect 81486 98758 81538 98810
rect 81538 98758 81540 98810
rect 81484 98756 81540 98758
rect 111996 98810 112052 98812
rect 111996 98758 111998 98810
rect 111998 98758 112050 98810
rect 112050 98758 112052 98810
rect 111996 98756 112052 98758
rect 112100 98810 112156 98812
rect 112100 98758 112102 98810
rect 112102 98758 112154 98810
rect 112154 98758 112156 98810
rect 112100 98756 112156 98758
rect 112204 98810 112260 98812
rect 112204 98758 112206 98810
rect 112206 98758 112258 98810
rect 112258 98758 112260 98810
rect 112204 98756 112260 98758
rect 118076 98140 118132 98196
rect 65916 98026 65972 98028
rect 65916 97974 65918 98026
rect 65918 97974 65970 98026
rect 65970 97974 65972 98026
rect 65916 97972 65972 97974
rect 66020 98026 66076 98028
rect 66020 97974 66022 98026
rect 66022 97974 66074 98026
rect 66074 97974 66076 98026
rect 66020 97972 66076 97974
rect 66124 98026 66180 98028
rect 66124 97974 66126 98026
rect 66126 97974 66178 98026
rect 66178 97974 66180 98026
rect 66124 97972 66180 97974
rect 96636 98026 96692 98028
rect 96636 97974 96638 98026
rect 96638 97974 96690 98026
rect 96690 97974 96692 98026
rect 96636 97972 96692 97974
rect 96740 98026 96796 98028
rect 96740 97974 96742 98026
rect 96742 97974 96794 98026
rect 96794 97974 96796 98026
rect 96740 97972 96796 97974
rect 96844 98026 96900 98028
rect 96844 97974 96846 98026
rect 96846 97974 96898 98026
rect 96898 97974 96900 98026
rect 96844 97972 96900 97974
rect 81276 97242 81332 97244
rect 81276 97190 81278 97242
rect 81278 97190 81330 97242
rect 81330 97190 81332 97242
rect 81276 97188 81332 97190
rect 81380 97242 81436 97244
rect 81380 97190 81382 97242
rect 81382 97190 81434 97242
rect 81434 97190 81436 97242
rect 81380 97188 81436 97190
rect 81484 97242 81540 97244
rect 81484 97190 81486 97242
rect 81486 97190 81538 97242
rect 81538 97190 81540 97242
rect 81484 97188 81540 97190
rect 111996 97242 112052 97244
rect 111996 97190 111998 97242
rect 111998 97190 112050 97242
rect 112050 97190 112052 97242
rect 111996 97188 112052 97190
rect 112100 97242 112156 97244
rect 112100 97190 112102 97242
rect 112102 97190 112154 97242
rect 112154 97190 112156 97242
rect 112100 97188 112156 97190
rect 112204 97242 112260 97244
rect 112204 97190 112206 97242
rect 112206 97190 112258 97242
rect 112258 97190 112260 97242
rect 112204 97188 112260 97190
rect 118076 96796 118132 96852
rect 65916 96458 65972 96460
rect 65916 96406 65918 96458
rect 65918 96406 65970 96458
rect 65970 96406 65972 96458
rect 65916 96404 65972 96406
rect 66020 96458 66076 96460
rect 66020 96406 66022 96458
rect 66022 96406 66074 96458
rect 66074 96406 66076 96458
rect 66020 96404 66076 96406
rect 66124 96458 66180 96460
rect 66124 96406 66126 96458
rect 66126 96406 66178 96458
rect 66178 96406 66180 96458
rect 66124 96404 66180 96406
rect 96636 96458 96692 96460
rect 96636 96406 96638 96458
rect 96638 96406 96690 96458
rect 96690 96406 96692 96458
rect 96636 96404 96692 96406
rect 96740 96458 96796 96460
rect 96740 96406 96742 96458
rect 96742 96406 96794 96458
rect 96794 96406 96796 96458
rect 96740 96404 96796 96406
rect 96844 96458 96900 96460
rect 96844 96406 96846 96458
rect 96846 96406 96898 96458
rect 96898 96406 96900 96458
rect 96844 96404 96900 96406
rect 81276 95674 81332 95676
rect 81276 95622 81278 95674
rect 81278 95622 81330 95674
rect 81330 95622 81332 95674
rect 81276 95620 81332 95622
rect 81380 95674 81436 95676
rect 81380 95622 81382 95674
rect 81382 95622 81434 95674
rect 81434 95622 81436 95674
rect 81380 95620 81436 95622
rect 81484 95674 81540 95676
rect 81484 95622 81486 95674
rect 81486 95622 81538 95674
rect 81538 95622 81540 95674
rect 81484 95620 81540 95622
rect 111996 95674 112052 95676
rect 111996 95622 111998 95674
rect 111998 95622 112050 95674
rect 112050 95622 112052 95674
rect 111996 95620 112052 95622
rect 112100 95674 112156 95676
rect 112100 95622 112102 95674
rect 112102 95622 112154 95674
rect 112154 95622 112156 95674
rect 112100 95620 112156 95622
rect 112204 95674 112260 95676
rect 112204 95622 112206 95674
rect 112206 95622 112258 95674
rect 112258 95622 112260 95674
rect 112204 95620 112260 95622
rect 118076 95452 118132 95508
rect 65916 94890 65972 94892
rect 65916 94838 65918 94890
rect 65918 94838 65970 94890
rect 65970 94838 65972 94890
rect 65916 94836 65972 94838
rect 66020 94890 66076 94892
rect 66020 94838 66022 94890
rect 66022 94838 66074 94890
rect 66074 94838 66076 94890
rect 66020 94836 66076 94838
rect 66124 94890 66180 94892
rect 66124 94838 66126 94890
rect 66126 94838 66178 94890
rect 66178 94838 66180 94890
rect 66124 94836 66180 94838
rect 96636 94890 96692 94892
rect 96636 94838 96638 94890
rect 96638 94838 96690 94890
rect 96690 94838 96692 94890
rect 96636 94836 96692 94838
rect 96740 94890 96796 94892
rect 96740 94838 96742 94890
rect 96742 94838 96794 94890
rect 96794 94838 96796 94890
rect 96740 94836 96796 94838
rect 96844 94890 96900 94892
rect 96844 94838 96846 94890
rect 96846 94838 96898 94890
rect 96898 94838 96900 94890
rect 96844 94836 96900 94838
rect 81276 94106 81332 94108
rect 81276 94054 81278 94106
rect 81278 94054 81330 94106
rect 81330 94054 81332 94106
rect 81276 94052 81332 94054
rect 81380 94106 81436 94108
rect 81380 94054 81382 94106
rect 81382 94054 81434 94106
rect 81434 94054 81436 94106
rect 81380 94052 81436 94054
rect 81484 94106 81540 94108
rect 81484 94054 81486 94106
rect 81486 94054 81538 94106
rect 81538 94054 81540 94106
rect 81484 94052 81540 94054
rect 111996 94106 112052 94108
rect 111996 94054 111998 94106
rect 111998 94054 112050 94106
rect 112050 94054 112052 94106
rect 111996 94052 112052 94054
rect 112100 94106 112156 94108
rect 112100 94054 112102 94106
rect 112102 94054 112154 94106
rect 112154 94054 112156 94106
rect 112100 94052 112156 94054
rect 112204 94106 112260 94108
rect 112204 94054 112206 94106
rect 112206 94054 112258 94106
rect 112258 94054 112260 94106
rect 112204 94052 112260 94054
rect 65916 93322 65972 93324
rect 65916 93270 65918 93322
rect 65918 93270 65970 93322
rect 65970 93270 65972 93322
rect 65916 93268 65972 93270
rect 66020 93322 66076 93324
rect 66020 93270 66022 93322
rect 66022 93270 66074 93322
rect 66074 93270 66076 93322
rect 66020 93268 66076 93270
rect 66124 93322 66180 93324
rect 66124 93270 66126 93322
rect 66126 93270 66178 93322
rect 66178 93270 66180 93322
rect 66124 93268 66180 93270
rect 96636 93322 96692 93324
rect 96636 93270 96638 93322
rect 96638 93270 96690 93322
rect 96690 93270 96692 93322
rect 96636 93268 96692 93270
rect 96740 93322 96796 93324
rect 96740 93270 96742 93322
rect 96742 93270 96794 93322
rect 96794 93270 96796 93322
rect 96740 93268 96796 93270
rect 96844 93322 96900 93324
rect 96844 93270 96846 93322
rect 96846 93270 96898 93322
rect 96898 93270 96900 93322
rect 96844 93268 96900 93270
rect 81276 92538 81332 92540
rect 81276 92486 81278 92538
rect 81278 92486 81330 92538
rect 81330 92486 81332 92538
rect 81276 92484 81332 92486
rect 81380 92538 81436 92540
rect 81380 92486 81382 92538
rect 81382 92486 81434 92538
rect 81434 92486 81436 92538
rect 81380 92484 81436 92486
rect 81484 92538 81540 92540
rect 81484 92486 81486 92538
rect 81486 92486 81538 92538
rect 81538 92486 81540 92538
rect 81484 92484 81540 92486
rect 111996 92538 112052 92540
rect 111996 92486 111998 92538
rect 111998 92486 112050 92538
rect 112050 92486 112052 92538
rect 111996 92484 112052 92486
rect 112100 92538 112156 92540
rect 112100 92486 112102 92538
rect 112102 92486 112154 92538
rect 112154 92486 112156 92538
rect 112100 92484 112156 92486
rect 112204 92538 112260 92540
rect 112204 92486 112206 92538
rect 112206 92486 112258 92538
rect 112258 92486 112260 92538
rect 112204 92484 112260 92486
rect 65916 91754 65972 91756
rect 65916 91702 65918 91754
rect 65918 91702 65970 91754
rect 65970 91702 65972 91754
rect 65916 91700 65972 91702
rect 66020 91754 66076 91756
rect 66020 91702 66022 91754
rect 66022 91702 66074 91754
rect 66074 91702 66076 91754
rect 66020 91700 66076 91702
rect 66124 91754 66180 91756
rect 66124 91702 66126 91754
rect 66126 91702 66178 91754
rect 66178 91702 66180 91754
rect 66124 91700 66180 91702
rect 96636 91754 96692 91756
rect 96636 91702 96638 91754
rect 96638 91702 96690 91754
rect 96690 91702 96692 91754
rect 96636 91700 96692 91702
rect 96740 91754 96796 91756
rect 96740 91702 96742 91754
rect 96742 91702 96794 91754
rect 96794 91702 96796 91754
rect 96740 91700 96796 91702
rect 96844 91754 96900 91756
rect 96844 91702 96846 91754
rect 96846 91702 96898 91754
rect 96898 91702 96900 91754
rect 96844 91700 96900 91702
rect 81276 90970 81332 90972
rect 81276 90918 81278 90970
rect 81278 90918 81330 90970
rect 81330 90918 81332 90970
rect 81276 90916 81332 90918
rect 81380 90970 81436 90972
rect 81380 90918 81382 90970
rect 81382 90918 81434 90970
rect 81434 90918 81436 90970
rect 81380 90916 81436 90918
rect 81484 90970 81540 90972
rect 81484 90918 81486 90970
rect 81486 90918 81538 90970
rect 81538 90918 81540 90970
rect 81484 90916 81540 90918
rect 111996 90970 112052 90972
rect 111996 90918 111998 90970
rect 111998 90918 112050 90970
rect 112050 90918 112052 90970
rect 111996 90916 112052 90918
rect 112100 90970 112156 90972
rect 112100 90918 112102 90970
rect 112102 90918 112154 90970
rect 112154 90918 112156 90970
rect 112100 90916 112156 90918
rect 112204 90970 112260 90972
rect 112204 90918 112206 90970
rect 112206 90918 112258 90970
rect 112258 90918 112260 90970
rect 112204 90916 112260 90918
rect 118076 90748 118132 90804
rect 65916 90186 65972 90188
rect 65916 90134 65918 90186
rect 65918 90134 65970 90186
rect 65970 90134 65972 90186
rect 65916 90132 65972 90134
rect 66020 90186 66076 90188
rect 66020 90134 66022 90186
rect 66022 90134 66074 90186
rect 66074 90134 66076 90186
rect 66020 90132 66076 90134
rect 66124 90186 66180 90188
rect 66124 90134 66126 90186
rect 66126 90134 66178 90186
rect 66178 90134 66180 90186
rect 66124 90132 66180 90134
rect 96636 90186 96692 90188
rect 96636 90134 96638 90186
rect 96638 90134 96690 90186
rect 96690 90134 96692 90186
rect 96636 90132 96692 90134
rect 96740 90186 96796 90188
rect 96740 90134 96742 90186
rect 96742 90134 96794 90186
rect 96794 90134 96796 90186
rect 96740 90132 96796 90134
rect 96844 90186 96900 90188
rect 96844 90134 96846 90186
rect 96846 90134 96898 90186
rect 96898 90134 96900 90186
rect 96844 90132 96900 90134
rect 81276 89402 81332 89404
rect 81276 89350 81278 89402
rect 81278 89350 81330 89402
rect 81330 89350 81332 89402
rect 81276 89348 81332 89350
rect 81380 89402 81436 89404
rect 81380 89350 81382 89402
rect 81382 89350 81434 89402
rect 81434 89350 81436 89402
rect 81380 89348 81436 89350
rect 81484 89402 81540 89404
rect 81484 89350 81486 89402
rect 81486 89350 81538 89402
rect 81538 89350 81540 89402
rect 81484 89348 81540 89350
rect 111996 89402 112052 89404
rect 111996 89350 111998 89402
rect 111998 89350 112050 89402
rect 112050 89350 112052 89402
rect 111996 89348 112052 89350
rect 112100 89402 112156 89404
rect 112100 89350 112102 89402
rect 112102 89350 112154 89402
rect 112154 89350 112156 89402
rect 112100 89348 112156 89350
rect 112204 89402 112260 89404
rect 112204 89350 112206 89402
rect 112206 89350 112258 89402
rect 112258 89350 112260 89402
rect 112204 89348 112260 89350
rect 65916 88618 65972 88620
rect 65916 88566 65918 88618
rect 65918 88566 65970 88618
rect 65970 88566 65972 88618
rect 65916 88564 65972 88566
rect 66020 88618 66076 88620
rect 66020 88566 66022 88618
rect 66022 88566 66074 88618
rect 66074 88566 66076 88618
rect 66020 88564 66076 88566
rect 66124 88618 66180 88620
rect 66124 88566 66126 88618
rect 66126 88566 66178 88618
rect 66178 88566 66180 88618
rect 66124 88564 66180 88566
rect 96636 88618 96692 88620
rect 96636 88566 96638 88618
rect 96638 88566 96690 88618
rect 96690 88566 96692 88618
rect 96636 88564 96692 88566
rect 96740 88618 96796 88620
rect 96740 88566 96742 88618
rect 96742 88566 96794 88618
rect 96794 88566 96796 88618
rect 96740 88564 96796 88566
rect 96844 88618 96900 88620
rect 96844 88566 96846 88618
rect 96846 88566 96898 88618
rect 96898 88566 96900 88618
rect 96844 88564 96900 88566
rect 118076 88114 118132 88116
rect 118076 88062 118078 88114
rect 118078 88062 118130 88114
rect 118130 88062 118132 88114
rect 118076 88060 118132 88062
rect 81276 87834 81332 87836
rect 81276 87782 81278 87834
rect 81278 87782 81330 87834
rect 81330 87782 81332 87834
rect 81276 87780 81332 87782
rect 81380 87834 81436 87836
rect 81380 87782 81382 87834
rect 81382 87782 81434 87834
rect 81434 87782 81436 87834
rect 81380 87780 81436 87782
rect 81484 87834 81540 87836
rect 81484 87782 81486 87834
rect 81486 87782 81538 87834
rect 81538 87782 81540 87834
rect 81484 87780 81540 87782
rect 111996 87834 112052 87836
rect 111996 87782 111998 87834
rect 111998 87782 112050 87834
rect 112050 87782 112052 87834
rect 111996 87780 112052 87782
rect 112100 87834 112156 87836
rect 112100 87782 112102 87834
rect 112102 87782 112154 87834
rect 112154 87782 112156 87834
rect 112100 87780 112156 87782
rect 112204 87834 112260 87836
rect 112204 87782 112206 87834
rect 112206 87782 112258 87834
rect 112258 87782 112260 87834
rect 112204 87780 112260 87782
rect 65916 87050 65972 87052
rect 65916 86998 65918 87050
rect 65918 86998 65970 87050
rect 65970 86998 65972 87050
rect 65916 86996 65972 86998
rect 66020 87050 66076 87052
rect 66020 86998 66022 87050
rect 66022 86998 66074 87050
rect 66074 86998 66076 87050
rect 66020 86996 66076 86998
rect 66124 87050 66180 87052
rect 66124 86998 66126 87050
rect 66126 86998 66178 87050
rect 66178 86998 66180 87050
rect 66124 86996 66180 86998
rect 96636 87050 96692 87052
rect 96636 86998 96638 87050
rect 96638 86998 96690 87050
rect 96690 86998 96692 87050
rect 96636 86996 96692 86998
rect 96740 87050 96796 87052
rect 96740 86998 96742 87050
rect 96742 86998 96794 87050
rect 96794 86998 96796 87050
rect 96740 86996 96796 86998
rect 96844 87050 96900 87052
rect 96844 86998 96846 87050
rect 96846 86998 96898 87050
rect 96898 86998 96900 87050
rect 96844 86996 96900 86998
rect 81276 86266 81332 86268
rect 81276 86214 81278 86266
rect 81278 86214 81330 86266
rect 81330 86214 81332 86266
rect 81276 86212 81332 86214
rect 81380 86266 81436 86268
rect 81380 86214 81382 86266
rect 81382 86214 81434 86266
rect 81434 86214 81436 86266
rect 81380 86212 81436 86214
rect 81484 86266 81540 86268
rect 81484 86214 81486 86266
rect 81486 86214 81538 86266
rect 81538 86214 81540 86266
rect 81484 86212 81540 86214
rect 111996 86266 112052 86268
rect 111996 86214 111998 86266
rect 111998 86214 112050 86266
rect 112050 86214 112052 86266
rect 111996 86212 112052 86214
rect 112100 86266 112156 86268
rect 112100 86214 112102 86266
rect 112102 86214 112154 86266
rect 112154 86214 112156 86266
rect 112100 86212 112156 86214
rect 112204 86266 112260 86268
rect 112204 86214 112206 86266
rect 112206 86214 112258 86266
rect 112258 86214 112260 86266
rect 112204 86212 112260 86214
rect 65916 85482 65972 85484
rect 65916 85430 65918 85482
rect 65918 85430 65970 85482
rect 65970 85430 65972 85482
rect 65916 85428 65972 85430
rect 66020 85482 66076 85484
rect 66020 85430 66022 85482
rect 66022 85430 66074 85482
rect 66074 85430 66076 85482
rect 66020 85428 66076 85430
rect 66124 85482 66180 85484
rect 66124 85430 66126 85482
rect 66126 85430 66178 85482
rect 66178 85430 66180 85482
rect 66124 85428 66180 85430
rect 96636 85482 96692 85484
rect 96636 85430 96638 85482
rect 96638 85430 96690 85482
rect 96690 85430 96692 85482
rect 96636 85428 96692 85430
rect 96740 85482 96796 85484
rect 96740 85430 96742 85482
rect 96742 85430 96794 85482
rect 96794 85430 96796 85482
rect 96740 85428 96796 85430
rect 96844 85482 96900 85484
rect 96844 85430 96846 85482
rect 96846 85430 96898 85482
rect 96898 85430 96900 85482
rect 96844 85428 96900 85430
rect 81276 84698 81332 84700
rect 81276 84646 81278 84698
rect 81278 84646 81330 84698
rect 81330 84646 81332 84698
rect 81276 84644 81332 84646
rect 81380 84698 81436 84700
rect 81380 84646 81382 84698
rect 81382 84646 81434 84698
rect 81434 84646 81436 84698
rect 81380 84644 81436 84646
rect 81484 84698 81540 84700
rect 81484 84646 81486 84698
rect 81486 84646 81538 84698
rect 81538 84646 81540 84698
rect 81484 84644 81540 84646
rect 111996 84698 112052 84700
rect 111996 84646 111998 84698
rect 111998 84646 112050 84698
rect 112050 84646 112052 84698
rect 111996 84644 112052 84646
rect 112100 84698 112156 84700
rect 112100 84646 112102 84698
rect 112102 84646 112154 84698
rect 112154 84646 112156 84698
rect 112100 84644 112156 84646
rect 112204 84698 112260 84700
rect 112204 84646 112206 84698
rect 112206 84646 112258 84698
rect 112258 84646 112260 84698
rect 112204 84644 112260 84646
rect 118076 84028 118132 84084
rect 65916 83914 65972 83916
rect 65916 83862 65918 83914
rect 65918 83862 65970 83914
rect 65970 83862 65972 83914
rect 65916 83860 65972 83862
rect 66020 83914 66076 83916
rect 66020 83862 66022 83914
rect 66022 83862 66074 83914
rect 66074 83862 66076 83914
rect 66020 83860 66076 83862
rect 66124 83914 66180 83916
rect 66124 83862 66126 83914
rect 66126 83862 66178 83914
rect 66178 83862 66180 83914
rect 66124 83860 66180 83862
rect 96636 83914 96692 83916
rect 96636 83862 96638 83914
rect 96638 83862 96690 83914
rect 96690 83862 96692 83914
rect 96636 83860 96692 83862
rect 96740 83914 96796 83916
rect 96740 83862 96742 83914
rect 96742 83862 96794 83914
rect 96794 83862 96796 83914
rect 96740 83860 96796 83862
rect 96844 83914 96900 83916
rect 96844 83862 96846 83914
rect 96846 83862 96898 83914
rect 96898 83862 96900 83914
rect 96844 83860 96900 83862
rect 81276 83130 81332 83132
rect 81276 83078 81278 83130
rect 81278 83078 81330 83130
rect 81330 83078 81332 83130
rect 81276 83076 81332 83078
rect 81380 83130 81436 83132
rect 81380 83078 81382 83130
rect 81382 83078 81434 83130
rect 81434 83078 81436 83130
rect 81380 83076 81436 83078
rect 81484 83130 81540 83132
rect 81484 83078 81486 83130
rect 81486 83078 81538 83130
rect 81538 83078 81540 83130
rect 81484 83076 81540 83078
rect 111996 83130 112052 83132
rect 111996 83078 111998 83130
rect 111998 83078 112050 83130
rect 112050 83078 112052 83130
rect 111996 83076 112052 83078
rect 112100 83130 112156 83132
rect 112100 83078 112102 83130
rect 112102 83078 112154 83130
rect 112154 83078 112156 83130
rect 112100 83076 112156 83078
rect 112204 83130 112260 83132
rect 112204 83078 112206 83130
rect 112206 83078 112258 83130
rect 112258 83078 112260 83130
rect 112204 83076 112260 83078
rect 65916 82346 65972 82348
rect 65916 82294 65918 82346
rect 65918 82294 65970 82346
rect 65970 82294 65972 82346
rect 65916 82292 65972 82294
rect 66020 82346 66076 82348
rect 66020 82294 66022 82346
rect 66022 82294 66074 82346
rect 66074 82294 66076 82346
rect 66020 82292 66076 82294
rect 66124 82346 66180 82348
rect 66124 82294 66126 82346
rect 66126 82294 66178 82346
rect 66178 82294 66180 82346
rect 66124 82292 66180 82294
rect 96636 82346 96692 82348
rect 96636 82294 96638 82346
rect 96638 82294 96690 82346
rect 96690 82294 96692 82346
rect 96636 82292 96692 82294
rect 96740 82346 96796 82348
rect 96740 82294 96742 82346
rect 96742 82294 96794 82346
rect 96794 82294 96796 82346
rect 96740 82292 96796 82294
rect 96844 82346 96900 82348
rect 96844 82294 96846 82346
rect 96846 82294 96898 82346
rect 96898 82294 96900 82346
rect 96844 82292 96900 82294
rect 118076 82012 118132 82068
rect 81276 81562 81332 81564
rect 81276 81510 81278 81562
rect 81278 81510 81330 81562
rect 81330 81510 81332 81562
rect 81276 81508 81332 81510
rect 81380 81562 81436 81564
rect 81380 81510 81382 81562
rect 81382 81510 81434 81562
rect 81434 81510 81436 81562
rect 81380 81508 81436 81510
rect 81484 81562 81540 81564
rect 81484 81510 81486 81562
rect 81486 81510 81538 81562
rect 81538 81510 81540 81562
rect 81484 81508 81540 81510
rect 111996 81562 112052 81564
rect 111996 81510 111998 81562
rect 111998 81510 112050 81562
rect 112050 81510 112052 81562
rect 111996 81508 112052 81510
rect 112100 81562 112156 81564
rect 112100 81510 112102 81562
rect 112102 81510 112154 81562
rect 112154 81510 112156 81562
rect 112100 81508 112156 81510
rect 112204 81562 112260 81564
rect 112204 81510 112206 81562
rect 112206 81510 112258 81562
rect 112258 81510 112260 81562
rect 112204 81508 112260 81510
rect 65916 80778 65972 80780
rect 65916 80726 65918 80778
rect 65918 80726 65970 80778
rect 65970 80726 65972 80778
rect 65916 80724 65972 80726
rect 66020 80778 66076 80780
rect 66020 80726 66022 80778
rect 66022 80726 66074 80778
rect 66074 80726 66076 80778
rect 66020 80724 66076 80726
rect 66124 80778 66180 80780
rect 66124 80726 66126 80778
rect 66126 80726 66178 80778
rect 66178 80726 66180 80778
rect 66124 80724 66180 80726
rect 96636 80778 96692 80780
rect 96636 80726 96638 80778
rect 96638 80726 96690 80778
rect 96690 80726 96692 80778
rect 96636 80724 96692 80726
rect 96740 80778 96796 80780
rect 96740 80726 96742 80778
rect 96742 80726 96794 80778
rect 96794 80726 96796 80778
rect 96740 80724 96796 80726
rect 96844 80778 96900 80780
rect 96844 80726 96846 80778
rect 96846 80726 96898 80778
rect 96898 80726 96900 80778
rect 96844 80724 96900 80726
rect 81276 79994 81332 79996
rect 81276 79942 81278 79994
rect 81278 79942 81330 79994
rect 81330 79942 81332 79994
rect 81276 79940 81332 79942
rect 81380 79994 81436 79996
rect 81380 79942 81382 79994
rect 81382 79942 81434 79994
rect 81434 79942 81436 79994
rect 81380 79940 81436 79942
rect 81484 79994 81540 79996
rect 81484 79942 81486 79994
rect 81486 79942 81538 79994
rect 81538 79942 81540 79994
rect 81484 79940 81540 79942
rect 111996 79994 112052 79996
rect 111996 79942 111998 79994
rect 111998 79942 112050 79994
rect 112050 79942 112052 79994
rect 111996 79940 112052 79942
rect 112100 79994 112156 79996
rect 112100 79942 112102 79994
rect 112102 79942 112154 79994
rect 112154 79942 112156 79994
rect 112100 79940 112156 79942
rect 112204 79994 112260 79996
rect 112204 79942 112206 79994
rect 112206 79942 112258 79994
rect 112258 79942 112260 79994
rect 112204 79940 112260 79942
rect 118076 79324 118132 79380
rect 65916 79210 65972 79212
rect 65916 79158 65918 79210
rect 65918 79158 65970 79210
rect 65970 79158 65972 79210
rect 65916 79156 65972 79158
rect 66020 79210 66076 79212
rect 66020 79158 66022 79210
rect 66022 79158 66074 79210
rect 66074 79158 66076 79210
rect 66020 79156 66076 79158
rect 66124 79210 66180 79212
rect 66124 79158 66126 79210
rect 66126 79158 66178 79210
rect 66178 79158 66180 79210
rect 66124 79156 66180 79158
rect 96636 79210 96692 79212
rect 96636 79158 96638 79210
rect 96638 79158 96690 79210
rect 96690 79158 96692 79210
rect 96636 79156 96692 79158
rect 96740 79210 96796 79212
rect 96740 79158 96742 79210
rect 96742 79158 96794 79210
rect 96794 79158 96796 79210
rect 96740 79156 96796 79158
rect 96844 79210 96900 79212
rect 96844 79158 96846 79210
rect 96846 79158 96898 79210
rect 96898 79158 96900 79210
rect 96844 79156 96900 79158
rect 81276 78426 81332 78428
rect 81276 78374 81278 78426
rect 81278 78374 81330 78426
rect 81330 78374 81332 78426
rect 81276 78372 81332 78374
rect 81380 78426 81436 78428
rect 81380 78374 81382 78426
rect 81382 78374 81434 78426
rect 81434 78374 81436 78426
rect 81380 78372 81436 78374
rect 81484 78426 81540 78428
rect 81484 78374 81486 78426
rect 81486 78374 81538 78426
rect 81538 78374 81540 78426
rect 81484 78372 81540 78374
rect 111996 78426 112052 78428
rect 111996 78374 111998 78426
rect 111998 78374 112050 78426
rect 112050 78374 112052 78426
rect 111996 78372 112052 78374
rect 112100 78426 112156 78428
rect 112100 78374 112102 78426
rect 112102 78374 112154 78426
rect 112154 78374 112156 78426
rect 112100 78372 112156 78374
rect 112204 78426 112260 78428
rect 112204 78374 112206 78426
rect 112206 78374 112258 78426
rect 112258 78374 112260 78426
rect 112204 78372 112260 78374
rect 65916 77642 65972 77644
rect 65916 77590 65918 77642
rect 65918 77590 65970 77642
rect 65970 77590 65972 77642
rect 65916 77588 65972 77590
rect 66020 77642 66076 77644
rect 66020 77590 66022 77642
rect 66022 77590 66074 77642
rect 66074 77590 66076 77642
rect 66020 77588 66076 77590
rect 66124 77642 66180 77644
rect 66124 77590 66126 77642
rect 66126 77590 66178 77642
rect 66178 77590 66180 77642
rect 66124 77588 66180 77590
rect 96636 77642 96692 77644
rect 96636 77590 96638 77642
rect 96638 77590 96690 77642
rect 96690 77590 96692 77642
rect 96636 77588 96692 77590
rect 96740 77642 96796 77644
rect 96740 77590 96742 77642
rect 96742 77590 96794 77642
rect 96794 77590 96796 77642
rect 96740 77588 96796 77590
rect 96844 77642 96900 77644
rect 96844 77590 96846 77642
rect 96846 77590 96898 77642
rect 96898 77590 96900 77642
rect 96844 77588 96900 77590
rect 81276 76858 81332 76860
rect 81276 76806 81278 76858
rect 81278 76806 81330 76858
rect 81330 76806 81332 76858
rect 81276 76804 81332 76806
rect 81380 76858 81436 76860
rect 81380 76806 81382 76858
rect 81382 76806 81434 76858
rect 81434 76806 81436 76858
rect 81380 76804 81436 76806
rect 81484 76858 81540 76860
rect 81484 76806 81486 76858
rect 81486 76806 81538 76858
rect 81538 76806 81540 76858
rect 81484 76804 81540 76806
rect 111996 76858 112052 76860
rect 111996 76806 111998 76858
rect 111998 76806 112050 76858
rect 112050 76806 112052 76858
rect 111996 76804 112052 76806
rect 112100 76858 112156 76860
rect 112100 76806 112102 76858
rect 112102 76806 112154 76858
rect 112154 76806 112156 76858
rect 112100 76804 112156 76806
rect 112204 76858 112260 76860
rect 112204 76806 112206 76858
rect 112206 76806 112258 76858
rect 112258 76806 112260 76858
rect 112204 76804 112260 76806
rect 118076 76636 118132 76692
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 96636 76074 96692 76076
rect 96636 76022 96638 76074
rect 96638 76022 96690 76074
rect 96690 76022 96692 76074
rect 96636 76020 96692 76022
rect 96740 76074 96796 76076
rect 96740 76022 96742 76074
rect 96742 76022 96794 76074
rect 96794 76022 96796 76074
rect 96740 76020 96796 76022
rect 96844 76074 96900 76076
rect 96844 76022 96846 76074
rect 96846 76022 96898 76074
rect 96898 76022 96900 76074
rect 96844 76020 96900 76022
rect 81276 75290 81332 75292
rect 81276 75238 81278 75290
rect 81278 75238 81330 75290
rect 81330 75238 81332 75290
rect 81276 75236 81332 75238
rect 81380 75290 81436 75292
rect 81380 75238 81382 75290
rect 81382 75238 81434 75290
rect 81434 75238 81436 75290
rect 81380 75236 81436 75238
rect 81484 75290 81540 75292
rect 81484 75238 81486 75290
rect 81486 75238 81538 75290
rect 81538 75238 81540 75290
rect 81484 75236 81540 75238
rect 111996 75290 112052 75292
rect 111996 75238 111998 75290
rect 111998 75238 112050 75290
rect 112050 75238 112052 75290
rect 111996 75236 112052 75238
rect 112100 75290 112156 75292
rect 112100 75238 112102 75290
rect 112102 75238 112154 75290
rect 112154 75238 112156 75290
rect 112100 75236 112156 75238
rect 112204 75290 112260 75292
rect 112204 75238 112206 75290
rect 112206 75238 112258 75290
rect 112258 75238 112260 75290
rect 112204 75236 112260 75238
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 96636 74506 96692 74508
rect 96636 74454 96638 74506
rect 96638 74454 96690 74506
rect 96690 74454 96692 74506
rect 96636 74452 96692 74454
rect 96740 74506 96796 74508
rect 96740 74454 96742 74506
rect 96742 74454 96794 74506
rect 96794 74454 96796 74506
rect 96740 74452 96796 74454
rect 96844 74506 96900 74508
rect 96844 74454 96846 74506
rect 96846 74454 96898 74506
rect 96898 74454 96900 74506
rect 96844 74452 96900 74454
rect 81276 73722 81332 73724
rect 81276 73670 81278 73722
rect 81278 73670 81330 73722
rect 81330 73670 81332 73722
rect 81276 73668 81332 73670
rect 81380 73722 81436 73724
rect 81380 73670 81382 73722
rect 81382 73670 81434 73722
rect 81434 73670 81436 73722
rect 81380 73668 81436 73670
rect 81484 73722 81540 73724
rect 81484 73670 81486 73722
rect 81486 73670 81538 73722
rect 81538 73670 81540 73722
rect 81484 73668 81540 73670
rect 111996 73722 112052 73724
rect 111996 73670 111998 73722
rect 111998 73670 112050 73722
rect 112050 73670 112052 73722
rect 111996 73668 112052 73670
rect 112100 73722 112156 73724
rect 112100 73670 112102 73722
rect 112102 73670 112154 73722
rect 112154 73670 112156 73722
rect 112100 73668 112156 73670
rect 112204 73722 112260 73724
rect 112204 73670 112206 73722
rect 112206 73670 112258 73722
rect 112258 73670 112260 73722
rect 112204 73668 112260 73670
rect 118076 73276 118132 73332
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 96636 72938 96692 72940
rect 96636 72886 96638 72938
rect 96638 72886 96690 72938
rect 96690 72886 96692 72938
rect 96636 72884 96692 72886
rect 96740 72938 96796 72940
rect 96740 72886 96742 72938
rect 96742 72886 96794 72938
rect 96794 72886 96796 72938
rect 96740 72884 96796 72886
rect 96844 72938 96900 72940
rect 96844 72886 96846 72938
rect 96846 72886 96898 72938
rect 96898 72886 96900 72938
rect 96844 72884 96900 72886
rect 81276 72154 81332 72156
rect 81276 72102 81278 72154
rect 81278 72102 81330 72154
rect 81330 72102 81332 72154
rect 81276 72100 81332 72102
rect 81380 72154 81436 72156
rect 81380 72102 81382 72154
rect 81382 72102 81434 72154
rect 81434 72102 81436 72154
rect 81380 72100 81436 72102
rect 81484 72154 81540 72156
rect 81484 72102 81486 72154
rect 81486 72102 81538 72154
rect 81538 72102 81540 72154
rect 81484 72100 81540 72102
rect 111996 72154 112052 72156
rect 111996 72102 111998 72154
rect 111998 72102 112050 72154
rect 112050 72102 112052 72154
rect 111996 72100 112052 72102
rect 112100 72154 112156 72156
rect 112100 72102 112102 72154
rect 112102 72102 112154 72154
rect 112154 72102 112156 72154
rect 112100 72100 112156 72102
rect 112204 72154 112260 72156
rect 112204 72102 112206 72154
rect 112206 72102 112258 72154
rect 112258 72102 112260 72154
rect 112204 72100 112260 72102
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 96636 71370 96692 71372
rect 96636 71318 96638 71370
rect 96638 71318 96690 71370
rect 96690 71318 96692 71370
rect 96636 71316 96692 71318
rect 96740 71370 96796 71372
rect 96740 71318 96742 71370
rect 96742 71318 96794 71370
rect 96794 71318 96796 71370
rect 96740 71316 96796 71318
rect 96844 71370 96900 71372
rect 96844 71318 96846 71370
rect 96846 71318 96898 71370
rect 96898 71318 96900 71370
rect 96844 71316 96900 71318
rect 81276 70586 81332 70588
rect 81276 70534 81278 70586
rect 81278 70534 81330 70586
rect 81330 70534 81332 70586
rect 81276 70532 81332 70534
rect 81380 70586 81436 70588
rect 81380 70534 81382 70586
rect 81382 70534 81434 70586
rect 81434 70534 81436 70586
rect 81380 70532 81436 70534
rect 81484 70586 81540 70588
rect 81484 70534 81486 70586
rect 81486 70534 81538 70586
rect 81538 70534 81540 70586
rect 81484 70532 81540 70534
rect 111996 70586 112052 70588
rect 111996 70534 111998 70586
rect 111998 70534 112050 70586
rect 112050 70534 112052 70586
rect 111996 70532 112052 70534
rect 112100 70586 112156 70588
rect 112100 70534 112102 70586
rect 112102 70534 112154 70586
rect 112154 70534 112156 70586
rect 112100 70532 112156 70534
rect 112204 70586 112260 70588
rect 112204 70534 112206 70586
rect 112206 70534 112258 70586
rect 112258 70534 112260 70586
rect 112204 70532 112260 70534
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 96636 69802 96692 69804
rect 96636 69750 96638 69802
rect 96638 69750 96690 69802
rect 96690 69750 96692 69802
rect 96636 69748 96692 69750
rect 96740 69802 96796 69804
rect 96740 69750 96742 69802
rect 96742 69750 96794 69802
rect 96794 69750 96796 69802
rect 96740 69748 96796 69750
rect 96844 69802 96900 69804
rect 96844 69750 96846 69802
rect 96846 69750 96898 69802
rect 96898 69750 96900 69802
rect 96844 69748 96900 69750
rect 118076 69298 118132 69300
rect 118076 69246 118078 69298
rect 118078 69246 118130 69298
rect 118130 69246 118132 69298
rect 118076 69244 118132 69246
rect 81276 69018 81332 69020
rect 81276 68966 81278 69018
rect 81278 68966 81330 69018
rect 81330 68966 81332 69018
rect 81276 68964 81332 68966
rect 81380 69018 81436 69020
rect 81380 68966 81382 69018
rect 81382 68966 81434 69018
rect 81434 68966 81436 69018
rect 81380 68964 81436 68966
rect 81484 69018 81540 69020
rect 81484 68966 81486 69018
rect 81486 68966 81538 69018
rect 81538 68966 81540 69018
rect 81484 68964 81540 68966
rect 111996 69018 112052 69020
rect 111996 68966 111998 69018
rect 111998 68966 112050 69018
rect 112050 68966 112052 69018
rect 111996 68964 112052 68966
rect 112100 69018 112156 69020
rect 112100 68966 112102 69018
rect 112102 68966 112154 69018
rect 112154 68966 112156 69018
rect 112100 68964 112156 68966
rect 112204 69018 112260 69020
rect 112204 68966 112206 69018
rect 112206 68966 112258 69018
rect 112258 68966 112260 69018
rect 112204 68964 112260 68966
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 96636 68234 96692 68236
rect 96636 68182 96638 68234
rect 96638 68182 96690 68234
rect 96690 68182 96692 68234
rect 96636 68180 96692 68182
rect 96740 68234 96796 68236
rect 96740 68182 96742 68234
rect 96742 68182 96794 68234
rect 96794 68182 96796 68234
rect 96740 68180 96796 68182
rect 96844 68234 96900 68236
rect 96844 68182 96846 68234
rect 96846 68182 96898 68234
rect 96898 68182 96900 68234
rect 96844 68180 96900 68182
rect 60620 67900 60676 67956
rect 118076 67900 118132 67956
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 20636 66780 20692 66836
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 4060 45276 4116 45332
rect 2604 45052 2660 45108
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 2268 40908 2324 40964
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 1820 40348 1876 40404
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 1820 39004 1876 39060
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 1820 36988 1876 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 1820 35644 1876 35700
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 1820 32956 1876 33012
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 1820 29596 1876 29652
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1820 25564 1876 25620
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 1820 22876 1876 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1820 20860 1876 20916
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 1820 18172 1876 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 1820 16828 1876 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 1820 10780 1876 10836
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 1820 7420 1876 7476
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 1820 6076 1876 6132
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 1820 4732 1876 4788
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 28 2268 84 2324
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 81276 67450 81332 67452
rect 81276 67398 81278 67450
rect 81278 67398 81330 67450
rect 81330 67398 81332 67450
rect 81276 67396 81332 67398
rect 81380 67450 81436 67452
rect 81380 67398 81382 67450
rect 81382 67398 81434 67450
rect 81434 67398 81436 67450
rect 81380 67396 81436 67398
rect 81484 67450 81540 67452
rect 81484 67398 81486 67450
rect 81486 67398 81538 67450
rect 81538 67398 81540 67450
rect 81484 67396 81540 67398
rect 111996 67450 112052 67452
rect 111996 67398 111998 67450
rect 111998 67398 112050 67450
rect 112050 67398 112052 67450
rect 111996 67396 112052 67398
rect 112100 67450 112156 67452
rect 112100 67398 112102 67450
rect 112102 67398 112154 67450
rect 112154 67398 112156 67450
rect 112100 67396 112156 67398
rect 112204 67450 112260 67452
rect 112204 67398 112206 67450
rect 112206 67398 112258 67450
rect 112258 67398 112260 67450
rect 112204 67396 112260 67398
rect 118076 67228 118132 67284
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 96636 66666 96692 66668
rect 96636 66614 96638 66666
rect 96638 66614 96690 66666
rect 96690 66614 96692 66666
rect 96636 66612 96692 66614
rect 96740 66666 96796 66668
rect 96740 66614 96742 66666
rect 96742 66614 96794 66666
rect 96794 66614 96796 66666
rect 96740 66612 96796 66614
rect 96844 66666 96900 66668
rect 96844 66614 96846 66666
rect 96846 66614 96898 66666
rect 96898 66614 96900 66666
rect 96844 66612 96900 66614
rect 81276 65882 81332 65884
rect 81276 65830 81278 65882
rect 81278 65830 81330 65882
rect 81330 65830 81332 65882
rect 81276 65828 81332 65830
rect 81380 65882 81436 65884
rect 81380 65830 81382 65882
rect 81382 65830 81434 65882
rect 81434 65830 81436 65882
rect 81380 65828 81436 65830
rect 81484 65882 81540 65884
rect 81484 65830 81486 65882
rect 81486 65830 81538 65882
rect 81538 65830 81540 65882
rect 81484 65828 81540 65830
rect 111996 65882 112052 65884
rect 111996 65830 111998 65882
rect 111998 65830 112050 65882
rect 112050 65830 112052 65882
rect 111996 65828 112052 65830
rect 112100 65882 112156 65884
rect 112100 65830 112102 65882
rect 112102 65830 112154 65882
rect 112154 65830 112156 65882
rect 112100 65828 112156 65830
rect 112204 65882 112260 65884
rect 112204 65830 112206 65882
rect 112206 65830 112258 65882
rect 112258 65830 112260 65882
rect 112204 65828 112260 65830
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 96636 65098 96692 65100
rect 96636 65046 96638 65098
rect 96638 65046 96690 65098
rect 96690 65046 96692 65098
rect 96636 65044 96692 65046
rect 96740 65098 96796 65100
rect 96740 65046 96742 65098
rect 96742 65046 96794 65098
rect 96794 65046 96796 65098
rect 96740 65044 96796 65046
rect 96844 65098 96900 65100
rect 96844 65046 96846 65098
rect 96846 65046 96898 65098
rect 96898 65046 96900 65098
rect 96844 65044 96900 65046
rect 81276 64314 81332 64316
rect 81276 64262 81278 64314
rect 81278 64262 81330 64314
rect 81330 64262 81332 64314
rect 81276 64260 81332 64262
rect 81380 64314 81436 64316
rect 81380 64262 81382 64314
rect 81382 64262 81434 64314
rect 81434 64262 81436 64314
rect 81380 64260 81436 64262
rect 81484 64314 81540 64316
rect 81484 64262 81486 64314
rect 81486 64262 81538 64314
rect 81538 64262 81540 64314
rect 81484 64260 81540 64262
rect 111996 64314 112052 64316
rect 111996 64262 111998 64314
rect 111998 64262 112050 64314
rect 112050 64262 112052 64314
rect 111996 64260 112052 64262
rect 112100 64314 112156 64316
rect 112100 64262 112102 64314
rect 112102 64262 112154 64314
rect 112154 64262 112156 64314
rect 112100 64260 112156 64262
rect 112204 64314 112260 64316
rect 112204 64262 112206 64314
rect 112206 64262 112258 64314
rect 112258 64262 112260 64314
rect 112204 64260 112260 64262
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 96636 63530 96692 63532
rect 96636 63478 96638 63530
rect 96638 63478 96690 63530
rect 96690 63478 96692 63530
rect 96636 63476 96692 63478
rect 96740 63530 96796 63532
rect 96740 63478 96742 63530
rect 96742 63478 96794 63530
rect 96794 63478 96796 63530
rect 96740 63476 96796 63478
rect 96844 63530 96900 63532
rect 96844 63478 96846 63530
rect 96846 63478 96898 63530
rect 96898 63478 96900 63530
rect 96844 63476 96900 63478
rect 81276 62746 81332 62748
rect 81276 62694 81278 62746
rect 81278 62694 81330 62746
rect 81330 62694 81332 62746
rect 81276 62692 81332 62694
rect 81380 62746 81436 62748
rect 81380 62694 81382 62746
rect 81382 62694 81434 62746
rect 81434 62694 81436 62746
rect 81380 62692 81436 62694
rect 81484 62746 81540 62748
rect 81484 62694 81486 62746
rect 81486 62694 81538 62746
rect 81538 62694 81540 62746
rect 81484 62692 81540 62694
rect 111996 62746 112052 62748
rect 111996 62694 111998 62746
rect 111998 62694 112050 62746
rect 112050 62694 112052 62746
rect 111996 62692 112052 62694
rect 112100 62746 112156 62748
rect 112100 62694 112102 62746
rect 112102 62694 112154 62746
rect 112154 62694 112156 62746
rect 112100 62692 112156 62694
rect 112204 62746 112260 62748
rect 112204 62694 112206 62746
rect 112206 62694 112258 62746
rect 112258 62694 112260 62746
rect 112204 62692 112260 62694
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 96636 61962 96692 61964
rect 96636 61910 96638 61962
rect 96638 61910 96690 61962
rect 96690 61910 96692 61962
rect 96636 61908 96692 61910
rect 96740 61962 96796 61964
rect 96740 61910 96742 61962
rect 96742 61910 96794 61962
rect 96794 61910 96796 61962
rect 96740 61908 96796 61910
rect 96844 61962 96900 61964
rect 96844 61910 96846 61962
rect 96846 61910 96898 61962
rect 96898 61910 96900 61962
rect 96844 61908 96900 61910
rect 81276 61178 81332 61180
rect 81276 61126 81278 61178
rect 81278 61126 81330 61178
rect 81330 61126 81332 61178
rect 81276 61124 81332 61126
rect 81380 61178 81436 61180
rect 81380 61126 81382 61178
rect 81382 61126 81434 61178
rect 81434 61126 81436 61178
rect 81380 61124 81436 61126
rect 81484 61178 81540 61180
rect 81484 61126 81486 61178
rect 81486 61126 81538 61178
rect 81538 61126 81540 61178
rect 81484 61124 81540 61126
rect 111996 61178 112052 61180
rect 111996 61126 111998 61178
rect 111998 61126 112050 61178
rect 112050 61126 112052 61178
rect 111996 61124 112052 61126
rect 112100 61178 112156 61180
rect 112100 61126 112102 61178
rect 112102 61126 112154 61178
rect 112154 61126 112156 61178
rect 112100 61124 112156 61126
rect 112204 61178 112260 61180
rect 112204 61126 112206 61178
rect 112206 61126 112258 61178
rect 112258 61126 112260 61178
rect 112204 61124 112260 61126
rect 118076 60508 118132 60564
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 96636 60394 96692 60396
rect 96636 60342 96638 60394
rect 96638 60342 96690 60394
rect 96690 60342 96692 60394
rect 96636 60340 96692 60342
rect 96740 60394 96796 60396
rect 96740 60342 96742 60394
rect 96742 60342 96794 60394
rect 96794 60342 96796 60394
rect 96740 60340 96796 60342
rect 96844 60394 96900 60396
rect 96844 60342 96846 60394
rect 96846 60342 96898 60394
rect 96898 60342 96900 60394
rect 96844 60340 96900 60342
rect 118076 59890 118132 59892
rect 118076 59838 118078 59890
rect 118078 59838 118130 59890
rect 118130 59838 118132 59890
rect 118076 59836 118132 59838
rect 81276 59610 81332 59612
rect 81276 59558 81278 59610
rect 81278 59558 81330 59610
rect 81330 59558 81332 59610
rect 81276 59556 81332 59558
rect 81380 59610 81436 59612
rect 81380 59558 81382 59610
rect 81382 59558 81434 59610
rect 81434 59558 81436 59610
rect 81380 59556 81436 59558
rect 81484 59610 81540 59612
rect 81484 59558 81486 59610
rect 81486 59558 81538 59610
rect 81538 59558 81540 59610
rect 81484 59556 81540 59558
rect 111996 59610 112052 59612
rect 111996 59558 111998 59610
rect 111998 59558 112050 59610
rect 112050 59558 112052 59610
rect 111996 59556 112052 59558
rect 112100 59610 112156 59612
rect 112100 59558 112102 59610
rect 112102 59558 112154 59610
rect 112154 59558 112156 59610
rect 112100 59556 112156 59558
rect 112204 59610 112260 59612
rect 112204 59558 112206 59610
rect 112206 59558 112258 59610
rect 112258 59558 112260 59610
rect 112204 59556 112260 59558
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 96636 58826 96692 58828
rect 96636 58774 96638 58826
rect 96638 58774 96690 58826
rect 96690 58774 96692 58826
rect 96636 58772 96692 58774
rect 96740 58826 96796 58828
rect 96740 58774 96742 58826
rect 96742 58774 96794 58826
rect 96794 58774 96796 58826
rect 96740 58772 96796 58774
rect 96844 58826 96900 58828
rect 96844 58774 96846 58826
rect 96846 58774 96898 58826
rect 96898 58774 96900 58826
rect 96844 58772 96900 58774
rect 118076 58492 118132 58548
rect 81276 58042 81332 58044
rect 81276 57990 81278 58042
rect 81278 57990 81330 58042
rect 81330 57990 81332 58042
rect 81276 57988 81332 57990
rect 81380 58042 81436 58044
rect 81380 57990 81382 58042
rect 81382 57990 81434 58042
rect 81434 57990 81436 58042
rect 81380 57988 81436 57990
rect 81484 58042 81540 58044
rect 81484 57990 81486 58042
rect 81486 57990 81538 58042
rect 81538 57990 81540 58042
rect 81484 57988 81540 57990
rect 111996 58042 112052 58044
rect 111996 57990 111998 58042
rect 111998 57990 112050 58042
rect 112050 57990 112052 58042
rect 111996 57988 112052 57990
rect 112100 58042 112156 58044
rect 112100 57990 112102 58042
rect 112102 57990 112154 58042
rect 112154 57990 112156 58042
rect 112100 57988 112156 57990
rect 112204 58042 112260 58044
rect 112204 57990 112206 58042
rect 112206 57990 112258 58042
rect 112258 57990 112260 58042
rect 112204 57988 112260 57990
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 96636 57258 96692 57260
rect 96636 57206 96638 57258
rect 96638 57206 96690 57258
rect 96690 57206 96692 57258
rect 96636 57204 96692 57206
rect 96740 57258 96796 57260
rect 96740 57206 96742 57258
rect 96742 57206 96794 57258
rect 96794 57206 96796 57258
rect 96740 57204 96796 57206
rect 96844 57258 96900 57260
rect 96844 57206 96846 57258
rect 96846 57206 96898 57258
rect 96898 57206 96900 57258
rect 96844 57204 96900 57206
rect 118076 57148 118132 57204
rect 81276 56474 81332 56476
rect 81276 56422 81278 56474
rect 81278 56422 81330 56474
rect 81330 56422 81332 56474
rect 81276 56420 81332 56422
rect 81380 56474 81436 56476
rect 81380 56422 81382 56474
rect 81382 56422 81434 56474
rect 81434 56422 81436 56474
rect 81380 56420 81436 56422
rect 81484 56474 81540 56476
rect 81484 56422 81486 56474
rect 81486 56422 81538 56474
rect 81538 56422 81540 56474
rect 81484 56420 81540 56422
rect 111996 56474 112052 56476
rect 111996 56422 111998 56474
rect 111998 56422 112050 56474
rect 112050 56422 112052 56474
rect 111996 56420 112052 56422
rect 112100 56474 112156 56476
rect 112100 56422 112102 56474
rect 112102 56422 112154 56474
rect 112154 56422 112156 56474
rect 112100 56420 112156 56422
rect 112204 56474 112260 56476
rect 112204 56422 112206 56474
rect 112206 56422 112258 56474
rect 112258 56422 112260 56474
rect 112204 56420 112260 56422
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 96636 55690 96692 55692
rect 96636 55638 96638 55690
rect 96638 55638 96690 55690
rect 96690 55638 96692 55690
rect 96636 55636 96692 55638
rect 96740 55690 96796 55692
rect 96740 55638 96742 55690
rect 96742 55638 96794 55690
rect 96794 55638 96796 55690
rect 96740 55636 96796 55638
rect 96844 55690 96900 55692
rect 96844 55638 96846 55690
rect 96846 55638 96898 55690
rect 96898 55638 96900 55690
rect 96844 55636 96900 55638
rect 81276 54906 81332 54908
rect 81276 54854 81278 54906
rect 81278 54854 81330 54906
rect 81330 54854 81332 54906
rect 81276 54852 81332 54854
rect 81380 54906 81436 54908
rect 81380 54854 81382 54906
rect 81382 54854 81434 54906
rect 81434 54854 81436 54906
rect 81380 54852 81436 54854
rect 81484 54906 81540 54908
rect 81484 54854 81486 54906
rect 81486 54854 81538 54906
rect 81538 54854 81540 54906
rect 81484 54852 81540 54854
rect 111996 54906 112052 54908
rect 111996 54854 111998 54906
rect 111998 54854 112050 54906
rect 112050 54854 112052 54906
rect 111996 54852 112052 54854
rect 112100 54906 112156 54908
rect 112100 54854 112102 54906
rect 112102 54854 112154 54906
rect 112154 54854 112156 54906
rect 112100 54852 112156 54854
rect 112204 54906 112260 54908
rect 112204 54854 112206 54906
rect 112206 54854 112258 54906
rect 112258 54854 112260 54906
rect 112204 54852 112260 54854
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 96636 54122 96692 54124
rect 96636 54070 96638 54122
rect 96638 54070 96690 54122
rect 96690 54070 96692 54122
rect 96636 54068 96692 54070
rect 96740 54122 96796 54124
rect 96740 54070 96742 54122
rect 96742 54070 96794 54122
rect 96794 54070 96796 54122
rect 96740 54068 96796 54070
rect 96844 54122 96900 54124
rect 96844 54070 96846 54122
rect 96846 54070 96898 54122
rect 96898 54070 96900 54122
rect 96844 54068 96900 54070
rect 81276 53338 81332 53340
rect 81276 53286 81278 53338
rect 81278 53286 81330 53338
rect 81330 53286 81332 53338
rect 81276 53284 81332 53286
rect 81380 53338 81436 53340
rect 81380 53286 81382 53338
rect 81382 53286 81434 53338
rect 81434 53286 81436 53338
rect 81380 53284 81436 53286
rect 81484 53338 81540 53340
rect 81484 53286 81486 53338
rect 81486 53286 81538 53338
rect 81538 53286 81540 53338
rect 81484 53284 81540 53286
rect 111996 53338 112052 53340
rect 111996 53286 111998 53338
rect 111998 53286 112050 53338
rect 112050 53286 112052 53338
rect 111996 53284 112052 53286
rect 112100 53338 112156 53340
rect 112100 53286 112102 53338
rect 112102 53286 112154 53338
rect 112154 53286 112156 53338
rect 112100 53284 112156 53286
rect 112204 53338 112260 53340
rect 112204 53286 112206 53338
rect 112206 53286 112258 53338
rect 112258 53286 112260 53338
rect 112204 53284 112260 53286
rect 118076 53228 118132 53284
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 96636 52554 96692 52556
rect 96636 52502 96638 52554
rect 96638 52502 96690 52554
rect 96690 52502 96692 52554
rect 96636 52500 96692 52502
rect 96740 52554 96796 52556
rect 96740 52502 96742 52554
rect 96742 52502 96794 52554
rect 96794 52502 96796 52554
rect 96740 52500 96796 52502
rect 96844 52554 96900 52556
rect 96844 52502 96846 52554
rect 96846 52502 96898 52554
rect 96898 52502 96900 52554
rect 96844 52500 96900 52502
rect 118076 52444 118132 52500
rect 81276 51770 81332 51772
rect 81276 51718 81278 51770
rect 81278 51718 81330 51770
rect 81330 51718 81332 51770
rect 81276 51716 81332 51718
rect 81380 51770 81436 51772
rect 81380 51718 81382 51770
rect 81382 51718 81434 51770
rect 81434 51718 81436 51770
rect 81380 51716 81436 51718
rect 81484 51770 81540 51772
rect 81484 51718 81486 51770
rect 81486 51718 81538 51770
rect 81538 51718 81540 51770
rect 81484 51716 81540 51718
rect 111996 51770 112052 51772
rect 111996 51718 111998 51770
rect 111998 51718 112050 51770
rect 112050 51718 112052 51770
rect 111996 51716 112052 51718
rect 112100 51770 112156 51772
rect 112100 51718 112102 51770
rect 112102 51718 112154 51770
rect 112154 51718 112156 51770
rect 112100 51716 112156 51718
rect 112204 51770 112260 51772
rect 112204 51718 112206 51770
rect 112206 51718 112258 51770
rect 112258 51718 112260 51770
rect 112204 51716 112260 51718
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 96636 50986 96692 50988
rect 96636 50934 96638 50986
rect 96638 50934 96690 50986
rect 96690 50934 96692 50986
rect 96636 50932 96692 50934
rect 96740 50986 96796 50988
rect 96740 50934 96742 50986
rect 96742 50934 96794 50986
rect 96794 50934 96796 50986
rect 96740 50932 96796 50934
rect 96844 50986 96900 50988
rect 96844 50934 96846 50986
rect 96846 50934 96898 50986
rect 96898 50934 96900 50986
rect 96844 50932 96900 50934
rect 81276 50202 81332 50204
rect 81276 50150 81278 50202
rect 81278 50150 81330 50202
rect 81330 50150 81332 50202
rect 81276 50148 81332 50150
rect 81380 50202 81436 50204
rect 81380 50150 81382 50202
rect 81382 50150 81434 50202
rect 81434 50150 81436 50202
rect 81380 50148 81436 50150
rect 81484 50202 81540 50204
rect 81484 50150 81486 50202
rect 81486 50150 81538 50202
rect 81538 50150 81540 50202
rect 81484 50148 81540 50150
rect 111996 50202 112052 50204
rect 111996 50150 111998 50202
rect 111998 50150 112050 50202
rect 112050 50150 112052 50202
rect 111996 50148 112052 50150
rect 112100 50202 112156 50204
rect 112100 50150 112102 50202
rect 112102 50150 112154 50202
rect 112154 50150 112156 50202
rect 112100 50148 112156 50150
rect 112204 50202 112260 50204
rect 112204 50150 112206 50202
rect 112206 50150 112258 50202
rect 112258 50150 112260 50202
rect 112204 50148 112260 50150
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 96636 49418 96692 49420
rect 96636 49366 96638 49418
rect 96638 49366 96690 49418
rect 96690 49366 96692 49418
rect 96636 49364 96692 49366
rect 96740 49418 96796 49420
rect 96740 49366 96742 49418
rect 96742 49366 96794 49418
rect 96794 49366 96796 49418
rect 96740 49364 96796 49366
rect 96844 49418 96900 49420
rect 96844 49366 96846 49418
rect 96846 49366 96898 49418
rect 96898 49366 96900 49418
rect 96844 49364 96900 49366
rect 81276 48634 81332 48636
rect 81276 48582 81278 48634
rect 81278 48582 81330 48634
rect 81330 48582 81332 48634
rect 81276 48580 81332 48582
rect 81380 48634 81436 48636
rect 81380 48582 81382 48634
rect 81382 48582 81434 48634
rect 81434 48582 81436 48634
rect 81380 48580 81436 48582
rect 81484 48634 81540 48636
rect 81484 48582 81486 48634
rect 81486 48582 81538 48634
rect 81538 48582 81540 48634
rect 81484 48580 81540 48582
rect 111996 48634 112052 48636
rect 111996 48582 111998 48634
rect 111998 48582 112050 48634
rect 112050 48582 112052 48634
rect 111996 48580 112052 48582
rect 112100 48634 112156 48636
rect 112100 48582 112102 48634
rect 112102 48582 112154 48634
rect 112154 48582 112156 48634
rect 112100 48580 112156 48582
rect 112204 48634 112260 48636
rect 112204 48582 112206 48634
rect 112206 48582 112258 48634
rect 112258 48582 112260 48634
rect 112204 48580 112260 48582
rect 59276 48076 59332 48132
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 96636 47850 96692 47852
rect 96636 47798 96638 47850
rect 96638 47798 96690 47850
rect 96690 47798 96692 47850
rect 96636 47796 96692 47798
rect 96740 47850 96796 47852
rect 96740 47798 96742 47850
rect 96742 47798 96794 47850
rect 96794 47798 96796 47850
rect 96740 47796 96796 47798
rect 96844 47850 96900 47852
rect 96844 47798 96846 47850
rect 96846 47798 96898 47850
rect 96898 47798 96900 47850
rect 96844 47796 96900 47798
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 81276 47066 81332 47068
rect 81276 47014 81278 47066
rect 81278 47014 81330 47066
rect 81330 47014 81332 47066
rect 81276 47012 81332 47014
rect 81380 47066 81436 47068
rect 81380 47014 81382 47066
rect 81382 47014 81434 47066
rect 81434 47014 81436 47066
rect 81380 47012 81436 47014
rect 81484 47066 81540 47068
rect 81484 47014 81486 47066
rect 81486 47014 81538 47066
rect 81538 47014 81540 47066
rect 81484 47012 81540 47014
rect 111996 47066 112052 47068
rect 111996 47014 111998 47066
rect 111998 47014 112050 47066
rect 112050 47014 112052 47066
rect 111996 47012 112052 47014
rect 112100 47066 112156 47068
rect 112100 47014 112102 47066
rect 112102 47014 112154 47066
rect 112154 47014 112156 47066
rect 112100 47012 112156 47014
rect 112204 47066 112260 47068
rect 112204 47014 112206 47066
rect 112206 47014 112258 47066
rect 112258 47014 112260 47066
rect 118076 47068 118132 47124
rect 112204 47012 112260 47014
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 96636 46282 96692 46284
rect 96636 46230 96638 46282
rect 96638 46230 96690 46282
rect 96690 46230 96692 46282
rect 96636 46228 96692 46230
rect 96740 46282 96796 46284
rect 96740 46230 96742 46282
rect 96742 46230 96794 46282
rect 96794 46230 96796 46282
rect 96740 46228 96796 46230
rect 96844 46282 96900 46284
rect 96844 46230 96846 46282
rect 96846 46230 96898 46282
rect 96898 46230 96900 46282
rect 96844 46228 96900 46230
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 81276 45498 81332 45500
rect 81276 45446 81278 45498
rect 81278 45446 81330 45498
rect 81330 45446 81332 45498
rect 81276 45444 81332 45446
rect 81380 45498 81436 45500
rect 81380 45446 81382 45498
rect 81382 45446 81434 45498
rect 81434 45446 81436 45498
rect 81380 45444 81436 45446
rect 81484 45498 81540 45500
rect 81484 45446 81486 45498
rect 81486 45446 81538 45498
rect 81538 45446 81540 45498
rect 81484 45444 81540 45446
rect 111996 45498 112052 45500
rect 111996 45446 111998 45498
rect 111998 45446 112050 45498
rect 112050 45446 112052 45498
rect 111996 45444 112052 45446
rect 112100 45498 112156 45500
rect 112100 45446 112102 45498
rect 112102 45446 112154 45498
rect 112154 45446 112156 45498
rect 112100 45444 112156 45446
rect 112204 45498 112260 45500
rect 112204 45446 112206 45498
rect 112206 45446 112258 45498
rect 112258 45446 112260 45498
rect 112204 45444 112260 45446
rect 118076 45052 118132 45108
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 96636 44714 96692 44716
rect 96636 44662 96638 44714
rect 96638 44662 96690 44714
rect 96690 44662 96692 44714
rect 96636 44660 96692 44662
rect 96740 44714 96796 44716
rect 96740 44662 96742 44714
rect 96742 44662 96794 44714
rect 96794 44662 96796 44714
rect 96740 44660 96796 44662
rect 96844 44714 96900 44716
rect 96844 44662 96846 44714
rect 96846 44662 96898 44714
rect 96898 44662 96900 44714
rect 96844 44660 96900 44662
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 81276 43930 81332 43932
rect 81276 43878 81278 43930
rect 81278 43878 81330 43930
rect 81330 43878 81332 43930
rect 81276 43876 81332 43878
rect 81380 43930 81436 43932
rect 81380 43878 81382 43930
rect 81382 43878 81434 43930
rect 81434 43878 81436 43930
rect 81380 43876 81436 43878
rect 81484 43930 81540 43932
rect 81484 43878 81486 43930
rect 81486 43878 81538 43930
rect 81538 43878 81540 43930
rect 81484 43876 81540 43878
rect 111996 43930 112052 43932
rect 111996 43878 111998 43930
rect 111998 43878 112050 43930
rect 112050 43878 112052 43930
rect 111996 43876 112052 43878
rect 112100 43930 112156 43932
rect 112100 43878 112102 43930
rect 112102 43878 112154 43930
rect 112154 43878 112156 43930
rect 112100 43876 112156 43878
rect 112204 43930 112260 43932
rect 112204 43878 112206 43930
rect 112206 43878 112258 43930
rect 112258 43878 112260 43930
rect 112204 43876 112260 43878
rect 118076 43708 118132 43764
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 96636 43146 96692 43148
rect 96636 43094 96638 43146
rect 96638 43094 96690 43146
rect 96690 43094 96692 43146
rect 96636 43092 96692 43094
rect 96740 43146 96796 43148
rect 96740 43094 96742 43146
rect 96742 43094 96794 43146
rect 96794 43094 96796 43146
rect 96740 43092 96796 43094
rect 96844 43146 96900 43148
rect 96844 43094 96846 43146
rect 96846 43094 96898 43146
rect 96898 43094 96900 43146
rect 96844 43092 96900 43094
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 81276 42362 81332 42364
rect 81276 42310 81278 42362
rect 81278 42310 81330 42362
rect 81330 42310 81332 42362
rect 81276 42308 81332 42310
rect 81380 42362 81436 42364
rect 81380 42310 81382 42362
rect 81382 42310 81434 42362
rect 81434 42310 81436 42362
rect 81380 42308 81436 42310
rect 81484 42362 81540 42364
rect 81484 42310 81486 42362
rect 81486 42310 81538 42362
rect 81538 42310 81540 42362
rect 81484 42308 81540 42310
rect 111996 42362 112052 42364
rect 111996 42310 111998 42362
rect 111998 42310 112050 42362
rect 112050 42310 112052 42362
rect 111996 42308 112052 42310
rect 112100 42362 112156 42364
rect 112100 42310 112102 42362
rect 112102 42310 112154 42362
rect 112154 42310 112156 42362
rect 112100 42308 112156 42310
rect 112204 42362 112260 42364
rect 112204 42310 112206 42362
rect 112206 42310 112258 42362
rect 112258 42310 112260 42362
rect 112204 42308 112260 42310
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 96636 41578 96692 41580
rect 96636 41526 96638 41578
rect 96638 41526 96690 41578
rect 96690 41526 96692 41578
rect 96636 41524 96692 41526
rect 96740 41578 96796 41580
rect 96740 41526 96742 41578
rect 96742 41526 96794 41578
rect 96794 41526 96796 41578
rect 96740 41524 96796 41526
rect 96844 41578 96900 41580
rect 96844 41526 96846 41578
rect 96846 41526 96898 41578
rect 96898 41526 96900 41578
rect 96844 41524 96900 41526
rect 59388 40962 59444 40964
rect 59388 40910 59390 40962
rect 59390 40910 59442 40962
rect 59442 40910 59444 40962
rect 59388 40908 59444 40910
rect 118076 41074 118132 41076
rect 118076 41022 118078 41074
rect 118078 41022 118130 41074
rect 118130 41022 118132 41074
rect 118076 41020 118132 41022
rect 59948 40908 60004 40964
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 81276 40794 81332 40796
rect 81276 40742 81278 40794
rect 81278 40742 81330 40794
rect 81330 40742 81332 40794
rect 81276 40740 81332 40742
rect 81380 40794 81436 40796
rect 81380 40742 81382 40794
rect 81382 40742 81434 40794
rect 81434 40742 81436 40794
rect 81380 40740 81436 40742
rect 81484 40794 81540 40796
rect 81484 40742 81486 40794
rect 81486 40742 81538 40794
rect 81538 40742 81540 40794
rect 81484 40740 81540 40742
rect 111996 40794 112052 40796
rect 111996 40742 111998 40794
rect 111998 40742 112050 40794
rect 112050 40742 112052 40794
rect 111996 40740 112052 40742
rect 112100 40794 112156 40796
rect 112100 40742 112102 40794
rect 112102 40742 112154 40794
rect 112154 40742 112156 40794
rect 112100 40740 112156 40742
rect 112204 40794 112260 40796
rect 112204 40742 112206 40794
rect 112206 40742 112258 40794
rect 112258 40742 112260 40794
rect 112204 40740 112260 40742
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 96636 40010 96692 40012
rect 96636 39958 96638 40010
rect 96638 39958 96690 40010
rect 96690 39958 96692 40010
rect 96636 39956 96692 39958
rect 96740 40010 96796 40012
rect 96740 39958 96742 40010
rect 96742 39958 96794 40010
rect 96794 39958 96796 40010
rect 96740 39956 96796 39958
rect 96844 40010 96900 40012
rect 96844 39958 96846 40010
rect 96846 39958 96898 40010
rect 96898 39958 96900 40010
rect 96844 39956 96900 39958
rect 81276 39226 81332 39228
rect 81276 39174 81278 39226
rect 81278 39174 81330 39226
rect 81330 39174 81332 39226
rect 81276 39172 81332 39174
rect 81380 39226 81436 39228
rect 81380 39174 81382 39226
rect 81382 39174 81434 39226
rect 81434 39174 81436 39226
rect 81380 39172 81436 39174
rect 81484 39226 81540 39228
rect 81484 39174 81486 39226
rect 81486 39174 81538 39226
rect 81538 39174 81540 39226
rect 81484 39172 81540 39174
rect 111996 39226 112052 39228
rect 111996 39174 111998 39226
rect 111998 39174 112050 39226
rect 112050 39174 112052 39226
rect 111996 39172 112052 39174
rect 112100 39226 112156 39228
rect 112100 39174 112102 39226
rect 112102 39174 112154 39226
rect 112154 39174 112156 39226
rect 112100 39172 112156 39174
rect 112204 39226 112260 39228
rect 112204 39174 112206 39226
rect 112206 39174 112258 39226
rect 112258 39174 112260 39226
rect 112204 39172 112260 39174
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 96636 38442 96692 38444
rect 96636 38390 96638 38442
rect 96638 38390 96690 38442
rect 96690 38390 96692 38442
rect 96636 38388 96692 38390
rect 96740 38442 96796 38444
rect 96740 38390 96742 38442
rect 96742 38390 96794 38442
rect 96794 38390 96796 38442
rect 96740 38388 96796 38390
rect 96844 38442 96900 38444
rect 96844 38390 96846 38442
rect 96846 38390 96898 38442
rect 96898 38390 96900 38442
rect 96844 38388 96900 38390
rect 118076 38332 118132 38388
rect 81276 37658 81332 37660
rect 81276 37606 81278 37658
rect 81278 37606 81330 37658
rect 81330 37606 81332 37658
rect 81276 37604 81332 37606
rect 81380 37658 81436 37660
rect 81380 37606 81382 37658
rect 81382 37606 81434 37658
rect 81434 37606 81436 37658
rect 81380 37604 81436 37606
rect 81484 37658 81540 37660
rect 81484 37606 81486 37658
rect 81486 37606 81538 37658
rect 81538 37606 81540 37658
rect 81484 37604 81540 37606
rect 111996 37658 112052 37660
rect 111996 37606 111998 37658
rect 111998 37606 112050 37658
rect 112050 37606 112052 37658
rect 111996 37604 112052 37606
rect 112100 37658 112156 37660
rect 112100 37606 112102 37658
rect 112102 37606 112154 37658
rect 112154 37606 112156 37658
rect 112100 37604 112156 37606
rect 112204 37658 112260 37660
rect 112204 37606 112206 37658
rect 112206 37606 112258 37658
rect 112258 37606 112260 37658
rect 112204 37604 112260 37606
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 96636 36874 96692 36876
rect 96636 36822 96638 36874
rect 96638 36822 96690 36874
rect 96690 36822 96692 36874
rect 96636 36820 96692 36822
rect 96740 36874 96796 36876
rect 96740 36822 96742 36874
rect 96742 36822 96794 36874
rect 96794 36822 96796 36874
rect 96740 36820 96796 36822
rect 96844 36874 96900 36876
rect 96844 36822 96846 36874
rect 96846 36822 96898 36874
rect 96898 36822 96900 36874
rect 96844 36820 96900 36822
rect 117740 36316 117796 36372
rect 81276 36090 81332 36092
rect 81276 36038 81278 36090
rect 81278 36038 81330 36090
rect 81330 36038 81332 36090
rect 81276 36036 81332 36038
rect 81380 36090 81436 36092
rect 81380 36038 81382 36090
rect 81382 36038 81434 36090
rect 81434 36038 81436 36090
rect 81380 36036 81436 36038
rect 81484 36090 81540 36092
rect 81484 36038 81486 36090
rect 81486 36038 81538 36090
rect 81538 36038 81540 36090
rect 81484 36036 81540 36038
rect 111996 36090 112052 36092
rect 111996 36038 111998 36090
rect 111998 36038 112050 36090
rect 112050 36038 112052 36090
rect 111996 36036 112052 36038
rect 112100 36090 112156 36092
rect 112100 36038 112102 36090
rect 112102 36038 112154 36090
rect 112154 36038 112156 36090
rect 112100 36036 112156 36038
rect 112204 36090 112260 36092
rect 112204 36038 112206 36090
rect 112206 36038 112258 36090
rect 112258 36038 112260 36090
rect 112204 36036 112260 36038
rect 60284 35532 60340 35588
rect 116284 35586 116340 35588
rect 116284 35534 116286 35586
rect 116286 35534 116338 35586
rect 116338 35534 116340 35586
rect 116284 35532 116340 35534
rect 116844 35532 116900 35588
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 96636 35306 96692 35308
rect 96636 35254 96638 35306
rect 96638 35254 96690 35306
rect 96690 35254 96692 35306
rect 96636 35252 96692 35254
rect 96740 35306 96796 35308
rect 96740 35254 96742 35306
rect 96742 35254 96794 35306
rect 96794 35254 96796 35306
rect 96740 35252 96796 35254
rect 96844 35306 96900 35308
rect 96844 35254 96846 35306
rect 96846 35254 96898 35306
rect 96898 35254 96900 35306
rect 96844 35252 96900 35254
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 81276 34522 81332 34524
rect 81276 34470 81278 34522
rect 81278 34470 81330 34522
rect 81330 34470 81332 34522
rect 81276 34468 81332 34470
rect 81380 34522 81436 34524
rect 81380 34470 81382 34522
rect 81382 34470 81434 34522
rect 81434 34470 81436 34522
rect 81380 34468 81436 34470
rect 81484 34522 81540 34524
rect 81484 34470 81486 34522
rect 81486 34470 81538 34522
rect 81538 34470 81540 34522
rect 81484 34468 81540 34470
rect 111996 34522 112052 34524
rect 111996 34470 111998 34522
rect 111998 34470 112050 34522
rect 112050 34470 112052 34522
rect 111996 34468 112052 34470
rect 112100 34522 112156 34524
rect 112100 34470 112102 34522
rect 112102 34470 112154 34522
rect 112154 34470 112156 34522
rect 112100 34468 112156 34470
rect 112204 34522 112260 34524
rect 112204 34470 112206 34522
rect 112206 34470 112258 34522
rect 112258 34470 112260 34522
rect 112204 34468 112260 34470
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 96636 33738 96692 33740
rect 96636 33686 96638 33738
rect 96638 33686 96690 33738
rect 96690 33686 96692 33738
rect 96636 33684 96692 33686
rect 96740 33738 96796 33740
rect 96740 33686 96742 33738
rect 96742 33686 96794 33738
rect 96794 33686 96796 33738
rect 96740 33684 96796 33686
rect 96844 33738 96900 33740
rect 96844 33686 96846 33738
rect 96846 33686 96898 33738
rect 96898 33686 96900 33738
rect 96844 33684 96900 33686
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 81276 32954 81332 32956
rect 81276 32902 81278 32954
rect 81278 32902 81330 32954
rect 81330 32902 81332 32954
rect 81276 32900 81332 32902
rect 81380 32954 81436 32956
rect 81380 32902 81382 32954
rect 81382 32902 81434 32954
rect 81434 32902 81436 32954
rect 81380 32900 81436 32902
rect 81484 32954 81540 32956
rect 81484 32902 81486 32954
rect 81486 32902 81538 32954
rect 81538 32902 81540 32954
rect 81484 32900 81540 32902
rect 111996 32954 112052 32956
rect 111996 32902 111998 32954
rect 111998 32902 112050 32954
rect 112050 32902 112052 32954
rect 111996 32900 112052 32902
rect 112100 32954 112156 32956
rect 112100 32902 112102 32954
rect 112102 32902 112154 32954
rect 112154 32902 112156 32954
rect 112100 32900 112156 32902
rect 112204 32954 112260 32956
rect 112204 32902 112206 32954
rect 112206 32902 112258 32954
rect 112258 32902 112260 32954
rect 112204 32900 112260 32902
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 96636 32170 96692 32172
rect 96636 32118 96638 32170
rect 96638 32118 96690 32170
rect 96690 32118 96692 32170
rect 96636 32116 96692 32118
rect 96740 32170 96796 32172
rect 96740 32118 96742 32170
rect 96742 32118 96794 32170
rect 96794 32118 96796 32170
rect 96740 32116 96796 32118
rect 96844 32170 96900 32172
rect 96844 32118 96846 32170
rect 96846 32118 96898 32170
rect 96898 32118 96900 32170
rect 96844 32116 96900 32118
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 81276 31386 81332 31388
rect 81276 31334 81278 31386
rect 81278 31334 81330 31386
rect 81330 31334 81332 31386
rect 81276 31332 81332 31334
rect 81380 31386 81436 31388
rect 81380 31334 81382 31386
rect 81382 31334 81434 31386
rect 81434 31334 81436 31386
rect 81380 31332 81436 31334
rect 81484 31386 81540 31388
rect 81484 31334 81486 31386
rect 81486 31334 81538 31386
rect 81538 31334 81540 31386
rect 81484 31332 81540 31334
rect 111996 31386 112052 31388
rect 111996 31334 111998 31386
rect 111998 31334 112050 31386
rect 112050 31334 112052 31386
rect 111996 31332 112052 31334
rect 112100 31386 112156 31388
rect 112100 31334 112102 31386
rect 112102 31334 112154 31386
rect 112154 31334 112156 31386
rect 112100 31332 112156 31334
rect 112204 31386 112260 31388
rect 112204 31334 112206 31386
rect 112206 31334 112258 31386
rect 112258 31334 112260 31386
rect 112204 31332 112260 31334
rect 118076 30940 118132 30996
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 96636 30602 96692 30604
rect 96636 30550 96638 30602
rect 96638 30550 96690 30602
rect 96690 30550 96692 30602
rect 96636 30548 96692 30550
rect 96740 30602 96796 30604
rect 96740 30550 96742 30602
rect 96742 30550 96794 30602
rect 96794 30550 96796 30602
rect 96740 30548 96796 30550
rect 96844 30602 96900 30604
rect 96844 30550 96846 30602
rect 96846 30550 96898 30602
rect 96898 30550 96900 30602
rect 96844 30548 96900 30550
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 81276 29818 81332 29820
rect 81276 29766 81278 29818
rect 81278 29766 81330 29818
rect 81330 29766 81332 29818
rect 81276 29764 81332 29766
rect 81380 29818 81436 29820
rect 81380 29766 81382 29818
rect 81382 29766 81434 29818
rect 81434 29766 81436 29818
rect 81380 29764 81436 29766
rect 81484 29818 81540 29820
rect 81484 29766 81486 29818
rect 81486 29766 81538 29818
rect 81538 29766 81540 29818
rect 81484 29764 81540 29766
rect 111996 29818 112052 29820
rect 111996 29766 111998 29818
rect 111998 29766 112050 29818
rect 112050 29766 112052 29818
rect 111996 29764 112052 29766
rect 112100 29818 112156 29820
rect 112100 29766 112102 29818
rect 112102 29766 112154 29818
rect 112154 29766 112156 29818
rect 112100 29764 112156 29766
rect 112204 29818 112260 29820
rect 112204 29766 112206 29818
rect 112206 29766 112258 29818
rect 112258 29766 112260 29818
rect 112204 29764 112260 29766
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 96636 29034 96692 29036
rect 96636 28982 96638 29034
rect 96638 28982 96690 29034
rect 96690 28982 96692 29034
rect 96636 28980 96692 28982
rect 96740 29034 96796 29036
rect 96740 28982 96742 29034
rect 96742 28982 96794 29034
rect 96794 28982 96796 29034
rect 96740 28980 96796 28982
rect 96844 29034 96900 29036
rect 96844 28982 96846 29034
rect 96846 28982 96898 29034
rect 96898 28982 96900 29034
rect 96844 28980 96900 28982
rect 118076 28924 118132 28980
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 81276 28250 81332 28252
rect 81276 28198 81278 28250
rect 81278 28198 81330 28250
rect 81330 28198 81332 28250
rect 81276 28196 81332 28198
rect 81380 28250 81436 28252
rect 81380 28198 81382 28250
rect 81382 28198 81434 28250
rect 81434 28198 81436 28250
rect 81380 28196 81436 28198
rect 81484 28250 81540 28252
rect 81484 28198 81486 28250
rect 81486 28198 81538 28250
rect 81538 28198 81540 28250
rect 81484 28196 81540 28198
rect 111996 28250 112052 28252
rect 111996 28198 111998 28250
rect 111998 28198 112050 28250
rect 112050 28198 112052 28250
rect 111996 28196 112052 28198
rect 112100 28250 112156 28252
rect 112100 28198 112102 28250
rect 112102 28198 112154 28250
rect 112154 28198 112156 28250
rect 112100 28196 112156 28198
rect 112204 28250 112260 28252
rect 112204 28198 112206 28250
rect 112206 28198 112258 28250
rect 112258 28198 112260 28250
rect 112204 28196 112260 28198
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 96636 27466 96692 27468
rect 96636 27414 96638 27466
rect 96638 27414 96690 27466
rect 96690 27414 96692 27466
rect 96636 27412 96692 27414
rect 96740 27466 96796 27468
rect 96740 27414 96742 27466
rect 96742 27414 96794 27466
rect 96794 27414 96796 27466
rect 96740 27412 96796 27414
rect 96844 27466 96900 27468
rect 96844 27414 96846 27466
rect 96846 27414 96898 27466
rect 96898 27414 96900 27466
rect 96844 27412 96900 27414
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 81276 26682 81332 26684
rect 81276 26630 81278 26682
rect 81278 26630 81330 26682
rect 81330 26630 81332 26682
rect 81276 26628 81332 26630
rect 81380 26682 81436 26684
rect 81380 26630 81382 26682
rect 81382 26630 81434 26682
rect 81434 26630 81436 26682
rect 81380 26628 81436 26630
rect 81484 26682 81540 26684
rect 81484 26630 81486 26682
rect 81486 26630 81538 26682
rect 81538 26630 81540 26682
rect 81484 26628 81540 26630
rect 111996 26682 112052 26684
rect 111996 26630 111998 26682
rect 111998 26630 112050 26682
rect 112050 26630 112052 26682
rect 111996 26628 112052 26630
rect 112100 26682 112156 26684
rect 112100 26630 112102 26682
rect 112102 26630 112154 26682
rect 112154 26630 112156 26682
rect 112100 26628 112156 26630
rect 112204 26682 112260 26684
rect 112204 26630 112206 26682
rect 112206 26630 112258 26682
rect 112258 26630 112260 26682
rect 112204 26628 112260 26630
rect 118076 26236 118132 26292
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 96636 25898 96692 25900
rect 96636 25846 96638 25898
rect 96638 25846 96690 25898
rect 96690 25846 96692 25898
rect 96636 25844 96692 25846
rect 96740 25898 96796 25900
rect 96740 25846 96742 25898
rect 96742 25846 96794 25898
rect 96794 25846 96796 25898
rect 96740 25844 96796 25846
rect 96844 25898 96900 25900
rect 96844 25846 96846 25898
rect 96846 25846 96898 25898
rect 96898 25846 96900 25898
rect 96844 25844 96900 25846
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 81276 25114 81332 25116
rect 81276 25062 81278 25114
rect 81278 25062 81330 25114
rect 81330 25062 81332 25114
rect 81276 25060 81332 25062
rect 81380 25114 81436 25116
rect 81380 25062 81382 25114
rect 81382 25062 81434 25114
rect 81434 25062 81436 25114
rect 81380 25060 81436 25062
rect 81484 25114 81540 25116
rect 81484 25062 81486 25114
rect 81486 25062 81538 25114
rect 81538 25062 81540 25114
rect 81484 25060 81540 25062
rect 111996 25114 112052 25116
rect 111996 25062 111998 25114
rect 111998 25062 112050 25114
rect 112050 25062 112052 25114
rect 111996 25060 112052 25062
rect 112100 25114 112156 25116
rect 112100 25062 112102 25114
rect 112102 25062 112154 25114
rect 112154 25062 112156 25114
rect 112100 25060 112156 25062
rect 112204 25114 112260 25116
rect 112204 25062 112206 25114
rect 112206 25062 112258 25114
rect 112258 25062 112260 25114
rect 112204 25060 112260 25062
rect 118076 24892 118132 24948
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 96636 24330 96692 24332
rect 96636 24278 96638 24330
rect 96638 24278 96690 24330
rect 96690 24278 96692 24330
rect 96636 24276 96692 24278
rect 96740 24330 96796 24332
rect 96740 24278 96742 24330
rect 96742 24278 96794 24330
rect 96794 24278 96796 24330
rect 96740 24276 96796 24278
rect 96844 24330 96900 24332
rect 96844 24278 96846 24330
rect 96846 24278 96898 24330
rect 96898 24278 96900 24330
rect 96844 24276 96900 24278
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 81276 23546 81332 23548
rect 81276 23494 81278 23546
rect 81278 23494 81330 23546
rect 81330 23494 81332 23546
rect 81276 23492 81332 23494
rect 81380 23546 81436 23548
rect 81380 23494 81382 23546
rect 81382 23494 81434 23546
rect 81434 23494 81436 23546
rect 81380 23492 81436 23494
rect 81484 23546 81540 23548
rect 81484 23494 81486 23546
rect 81486 23494 81538 23546
rect 81538 23494 81540 23546
rect 81484 23492 81540 23494
rect 111996 23546 112052 23548
rect 111996 23494 111998 23546
rect 111998 23494 112050 23546
rect 112050 23494 112052 23546
rect 111996 23492 112052 23494
rect 112100 23546 112156 23548
rect 112100 23494 112102 23546
rect 112102 23494 112154 23546
rect 112154 23494 112156 23546
rect 112100 23492 112156 23494
rect 112204 23546 112260 23548
rect 112204 23494 112206 23546
rect 112206 23494 112258 23546
rect 112258 23494 112260 23546
rect 112204 23492 112260 23494
rect 118076 22876 118132 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 96636 22762 96692 22764
rect 96636 22710 96638 22762
rect 96638 22710 96690 22762
rect 96690 22710 96692 22762
rect 96636 22708 96692 22710
rect 96740 22762 96796 22764
rect 96740 22710 96742 22762
rect 96742 22710 96794 22762
rect 96794 22710 96796 22762
rect 96740 22708 96796 22710
rect 96844 22762 96900 22764
rect 96844 22710 96846 22762
rect 96846 22710 96898 22762
rect 96898 22710 96900 22762
rect 96844 22708 96900 22710
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 81276 21978 81332 21980
rect 81276 21926 81278 21978
rect 81278 21926 81330 21978
rect 81330 21926 81332 21978
rect 81276 21924 81332 21926
rect 81380 21978 81436 21980
rect 81380 21926 81382 21978
rect 81382 21926 81434 21978
rect 81434 21926 81436 21978
rect 81380 21924 81436 21926
rect 81484 21978 81540 21980
rect 81484 21926 81486 21978
rect 81486 21926 81538 21978
rect 81538 21926 81540 21978
rect 81484 21924 81540 21926
rect 111996 21978 112052 21980
rect 111996 21926 111998 21978
rect 111998 21926 112050 21978
rect 112050 21926 112052 21978
rect 111996 21924 112052 21926
rect 112100 21978 112156 21980
rect 112100 21926 112102 21978
rect 112102 21926 112154 21978
rect 112154 21926 112156 21978
rect 112100 21924 112156 21926
rect 112204 21978 112260 21980
rect 112204 21926 112206 21978
rect 112206 21926 112258 21978
rect 112258 21926 112260 21978
rect 112204 21924 112260 21926
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 96636 21194 96692 21196
rect 96636 21142 96638 21194
rect 96638 21142 96690 21194
rect 96690 21142 96692 21194
rect 96636 21140 96692 21142
rect 96740 21194 96796 21196
rect 96740 21142 96742 21194
rect 96742 21142 96794 21194
rect 96794 21142 96796 21194
rect 96740 21140 96796 21142
rect 96844 21194 96900 21196
rect 96844 21142 96846 21194
rect 96846 21142 96898 21194
rect 96898 21142 96900 21194
rect 96844 21140 96900 21142
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 81276 20410 81332 20412
rect 81276 20358 81278 20410
rect 81278 20358 81330 20410
rect 81330 20358 81332 20410
rect 81276 20356 81332 20358
rect 81380 20410 81436 20412
rect 81380 20358 81382 20410
rect 81382 20358 81434 20410
rect 81434 20358 81436 20410
rect 81380 20356 81436 20358
rect 81484 20410 81540 20412
rect 81484 20358 81486 20410
rect 81486 20358 81538 20410
rect 81538 20358 81540 20410
rect 81484 20356 81540 20358
rect 111996 20410 112052 20412
rect 111996 20358 111998 20410
rect 111998 20358 112050 20410
rect 112050 20358 112052 20410
rect 111996 20356 112052 20358
rect 112100 20410 112156 20412
rect 112100 20358 112102 20410
rect 112102 20358 112154 20410
rect 112154 20358 112156 20410
rect 112100 20356 112156 20358
rect 112204 20410 112260 20412
rect 112204 20358 112206 20410
rect 112206 20358 112258 20410
rect 112258 20358 112260 20410
rect 112204 20356 112260 20358
rect 118076 20188 118132 20244
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 96636 19626 96692 19628
rect 96636 19574 96638 19626
rect 96638 19574 96690 19626
rect 96690 19574 96692 19626
rect 96636 19572 96692 19574
rect 96740 19626 96796 19628
rect 96740 19574 96742 19626
rect 96742 19574 96794 19626
rect 96794 19574 96796 19626
rect 96740 19572 96796 19574
rect 96844 19626 96900 19628
rect 96844 19574 96846 19626
rect 96846 19574 96898 19626
rect 96898 19574 96900 19626
rect 96844 19572 96900 19574
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 81276 18842 81332 18844
rect 81276 18790 81278 18842
rect 81278 18790 81330 18842
rect 81330 18790 81332 18842
rect 81276 18788 81332 18790
rect 81380 18842 81436 18844
rect 81380 18790 81382 18842
rect 81382 18790 81434 18842
rect 81434 18790 81436 18842
rect 81380 18788 81436 18790
rect 81484 18842 81540 18844
rect 81484 18790 81486 18842
rect 81486 18790 81538 18842
rect 81538 18790 81540 18842
rect 81484 18788 81540 18790
rect 111996 18842 112052 18844
rect 111996 18790 111998 18842
rect 111998 18790 112050 18842
rect 112050 18790 112052 18842
rect 111996 18788 112052 18790
rect 112100 18842 112156 18844
rect 112100 18790 112102 18842
rect 112102 18790 112154 18842
rect 112154 18790 112156 18842
rect 112100 18788 112156 18790
rect 112204 18842 112260 18844
rect 112204 18790 112206 18842
rect 112206 18790 112258 18842
rect 112258 18790 112260 18842
rect 112204 18788 112260 18790
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 96636 18058 96692 18060
rect 96636 18006 96638 18058
rect 96638 18006 96690 18058
rect 96690 18006 96692 18058
rect 96636 18004 96692 18006
rect 96740 18058 96796 18060
rect 96740 18006 96742 18058
rect 96742 18006 96794 18058
rect 96794 18006 96796 18058
rect 96740 18004 96796 18006
rect 96844 18058 96900 18060
rect 96844 18006 96846 18058
rect 96846 18006 96898 18058
rect 96898 18006 96900 18058
rect 96844 18004 96900 18006
rect 118076 17554 118132 17556
rect 118076 17502 118078 17554
rect 118078 17502 118130 17554
rect 118130 17502 118132 17554
rect 118076 17500 118132 17502
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 81276 17274 81332 17276
rect 81276 17222 81278 17274
rect 81278 17222 81330 17274
rect 81330 17222 81332 17274
rect 81276 17220 81332 17222
rect 81380 17274 81436 17276
rect 81380 17222 81382 17274
rect 81382 17222 81434 17274
rect 81434 17222 81436 17274
rect 81380 17220 81436 17222
rect 81484 17274 81540 17276
rect 81484 17222 81486 17274
rect 81486 17222 81538 17274
rect 81538 17222 81540 17274
rect 81484 17220 81540 17222
rect 111996 17274 112052 17276
rect 111996 17222 111998 17274
rect 111998 17222 112050 17274
rect 112050 17222 112052 17274
rect 111996 17220 112052 17222
rect 112100 17274 112156 17276
rect 112100 17222 112102 17274
rect 112102 17222 112154 17274
rect 112154 17222 112156 17274
rect 112100 17220 112156 17222
rect 112204 17274 112260 17276
rect 112204 17222 112206 17274
rect 112206 17222 112258 17274
rect 112258 17222 112260 17274
rect 112204 17220 112260 17222
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 96636 16490 96692 16492
rect 96636 16438 96638 16490
rect 96638 16438 96690 16490
rect 96690 16438 96692 16490
rect 96636 16436 96692 16438
rect 96740 16490 96796 16492
rect 96740 16438 96742 16490
rect 96742 16438 96794 16490
rect 96794 16438 96796 16490
rect 96740 16436 96796 16438
rect 96844 16490 96900 16492
rect 96844 16438 96846 16490
rect 96846 16438 96898 16490
rect 96898 16438 96900 16490
rect 96844 16436 96900 16438
rect 118076 16156 118132 16212
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 81276 15706 81332 15708
rect 81276 15654 81278 15706
rect 81278 15654 81330 15706
rect 81330 15654 81332 15706
rect 81276 15652 81332 15654
rect 81380 15706 81436 15708
rect 81380 15654 81382 15706
rect 81382 15654 81434 15706
rect 81434 15654 81436 15706
rect 81380 15652 81436 15654
rect 81484 15706 81540 15708
rect 81484 15654 81486 15706
rect 81486 15654 81538 15706
rect 81538 15654 81540 15706
rect 81484 15652 81540 15654
rect 111996 15706 112052 15708
rect 111996 15654 111998 15706
rect 111998 15654 112050 15706
rect 112050 15654 112052 15706
rect 111996 15652 112052 15654
rect 112100 15706 112156 15708
rect 112100 15654 112102 15706
rect 112102 15654 112154 15706
rect 112154 15654 112156 15706
rect 112100 15652 112156 15654
rect 112204 15706 112260 15708
rect 112204 15654 112206 15706
rect 112206 15654 112258 15706
rect 112258 15654 112260 15706
rect 112204 15652 112260 15654
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 96636 14922 96692 14924
rect 96636 14870 96638 14922
rect 96638 14870 96690 14922
rect 96690 14870 96692 14922
rect 96636 14868 96692 14870
rect 96740 14922 96796 14924
rect 96740 14870 96742 14922
rect 96742 14870 96794 14922
rect 96794 14870 96796 14922
rect 96740 14868 96796 14870
rect 96844 14922 96900 14924
rect 96844 14870 96846 14922
rect 96846 14870 96898 14922
rect 96898 14870 96900 14922
rect 96844 14868 96900 14870
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 81276 14138 81332 14140
rect 81276 14086 81278 14138
rect 81278 14086 81330 14138
rect 81330 14086 81332 14138
rect 81276 14084 81332 14086
rect 81380 14138 81436 14140
rect 81380 14086 81382 14138
rect 81382 14086 81434 14138
rect 81434 14086 81436 14138
rect 81380 14084 81436 14086
rect 81484 14138 81540 14140
rect 81484 14086 81486 14138
rect 81486 14086 81538 14138
rect 81538 14086 81540 14138
rect 81484 14084 81540 14086
rect 111996 14138 112052 14140
rect 111996 14086 111998 14138
rect 111998 14086 112050 14138
rect 112050 14086 112052 14138
rect 111996 14084 112052 14086
rect 112100 14138 112156 14140
rect 112100 14086 112102 14138
rect 112102 14086 112154 14138
rect 112154 14086 112156 14138
rect 112100 14084 112156 14086
rect 112204 14138 112260 14140
rect 112204 14086 112206 14138
rect 112206 14086 112258 14138
rect 112258 14086 112260 14138
rect 118076 14140 118132 14196
rect 112204 14084 112260 14086
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 96636 13354 96692 13356
rect 96636 13302 96638 13354
rect 96638 13302 96690 13354
rect 96690 13302 96692 13354
rect 96636 13300 96692 13302
rect 96740 13354 96796 13356
rect 96740 13302 96742 13354
rect 96742 13302 96794 13354
rect 96794 13302 96796 13354
rect 96740 13300 96796 13302
rect 96844 13354 96900 13356
rect 96844 13302 96846 13354
rect 96846 13302 96898 13354
rect 96898 13302 96900 13354
rect 96844 13300 96900 13302
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 81276 12570 81332 12572
rect 81276 12518 81278 12570
rect 81278 12518 81330 12570
rect 81330 12518 81332 12570
rect 81276 12516 81332 12518
rect 81380 12570 81436 12572
rect 81380 12518 81382 12570
rect 81382 12518 81434 12570
rect 81434 12518 81436 12570
rect 81380 12516 81436 12518
rect 81484 12570 81540 12572
rect 81484 12518 81486 12570
rect 81486 12518 81538 12570
rect 81538 12518 81540 12570
rect 81484 12516 81540 12518
rect 111996 12570 112052 12572
rect 111996 12518 111998 12570
rect 111998 12518 112050 12570
rect 112050 12518 112052 12570
rect 111996 12516 112052 12518
rect 112100 12570 112156 12572
rect 112100 12518 112102 12570
rect 112102 12518 112154 12570
rect 112154 12518 112156 12570
rect 112100 12516 112156 12518
rect 112204 12570 112260 12572
rect 112204 12518 112206 12570
rect 112206 12518 112258 12570
rect 112258 12518 112260 12570
rect 112204 12516 112260 12518
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 96636 11786 96692 11788
rect 96636 11734 96638 11786
rect 96638 11734 96690 11786
rect 96690 11734 96692 11786
rect 96636 11732 96692 11734
rect 96740 11786 96796 11788
rect 96740 11734 96742 11786
rect 96742 11734 96794 11786
rect 96794 11734 96796 11786
rect 96740 11732 96796 11734
rect 96844 11786 96900 11788
rect 96844 11734 96846 11786
rect 96846 11734 96898 11786
rect 96898 11734 96900 11786
rect 96844 11732 96900 11734
rect 118076 11452 118132 11508
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 81276 11002 81332 11004
rect 81276 10950 81278 11002
rect 81278 10950 81330 11002
rect 81330 10950 81332 11002
rect 81276 10948 81332 10950
rect 81380 11002 81436 11004
rect 81380 10950 81382 11002
rect 81382 10950 81434 11002
rect 81434 10950 81436 11002
rect 81380 10948 81436 10950
rect 81484 11002 81540 11004
rect 81484 10950 81486 11002
rect 81486 10950 81538 11002
rect 81538 10950 81540 11002
rect 81484 10948 81540 10950
rect 111996 11002 112052 11004
rect 111996 10950 111998 11002
rect 111998 10950 112050 11002
rect 112050 10950 112052 11002
rect 111996 10948 112052 10950
rect 112100 11002 112156 11004
rect 112100 10950 112102 11002
rect 112102 10950 112154 11002
rect 112154 10950 112156 11002
rect 112100 10948 112156 10950
rect 112204 11002 112260 11004
rect 112204 10950 112206 11002
rect 112206 10950 112258 11002
rect 112258 10950 112260 11002
rect 112204 10948 112260 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 96636 10218 96692 10220
rect 96636 10166 96638 10218
rect 96638 10166 96690 10218
rect 96690 10166 96692 10218
rect 96636 10164 96692 10166
rect 96740 10218 96796 10220
rect 96740 10166 96742 10218
rect 96742 10166 96794 10218
rect 96794 10166 96796 10218
rect 96740 10164 96796 10166
rect 96844 10218 96900 10220
rect 96844 10166 96846 10218
rect 96846 10166 96898 10218
rect 96898 10166 96900 10218
rect 96844 10164 96900 10166
rect 118076 10108 118132 10164
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 81276 9434 81332 9436
rect 81276 9382 81278 9434
rect 81278 9382 81330 9434
rect 81330 9382 81332 9434
rect 81276 9380 81332 9382
rect 81380 9434 81436 9436
rect 81380 9382 81382 9434
rect 81382 9382 81434 9434
rect 81434 9382 81436 9434
rect 81380 9380 81436 9382
rect 81484 9434 81540 9436
rect 81484 9382 81486 9434
rect 81486 9382 81538 9434
rect 81538 9382 81540 9434
rect 81484 9380 81540 9382
rect 111996 9434 112052 9436
rect 111996 9382 111998 9434
rect 111998 9382 112050 9434
rect 112050 9382 112052 9434
rect 111996 9380 112052 9382
rect 112100 9434 112156 9436
rect 112100 9382 112102 9434
rect 112102 9382 112154 9434
rect 112154 9382 112156 9434
rect 112100 9380 112156 9382
rect 112204 9434 112260 9436
rect 112204 9382 112206 9434
rect 112206 9382 112258 9434
rect 112258 9382 112260 9434
rect 112204 9380 112260 9382
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 96636 8650 96692 8652
rect 96636 8598 96638 8650
rect 96638 8598 96690 8650
rect 96690 8598 96692 8650
rect 96636 8596 96692 8598
rect 96740 8650 96796 8652
rect 96740 8598 96742 8650
rect 96742 8598 96794 8650
rect 96794 8598 96796 8650
rect 96740 8596 96796 8598
rect 96844 8650 96900 8652
rect 96844 8598 96846 8650
rect 96846 8598 96898 8650
rect 96898 8598 96900 8650
rect 96844 8596 96900 8598
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 81276 7866 81332 7868
rect 81276 7814 81278 7866
rect 81278 7814 81330 7866
rect 81330 7814 81332 7866
rect 81276 7812 81332 7814
rect 81380 7866 81436 7868
rect 81380 7814 81382 7866
rect 81382 7814 81434 7866
rect 81434 7814 81436 7866
rect 81380 7812 81436 7814
rect 81484 7866 81540 7868
rect 81484 7814 81486 7866
rect 81486 7814 81538 7866
rect 81538 7814 81540 7866
rect 81484 7812 81540 7814
rect 111996 7866 112052 7868
rect 111996 7814 111998 7866
rect 111998 7814 112050 7866
rect 112050 7814 112052 7866
rect 111996 7812 112052 7814
rect 112100 7866 112156 7868
rect 112100 7814 112102 7866
rect 112102 7814 112154 7866
rect 112154 7814 112156 7866
rect 112100 7812 112156 7814
rect 112204 7866 112260 7868
rect 112204 7814 112206 7866
rect 112206 7814 112258 7866
rect 112258 7814 112260 7866
rect 112204 7812 112260 7814
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 96636 7082 96692 7084
rect 96636 7030 96638 7082
rect 96638 7030 96690 7082
rect 96690 7030 96692 7082
rect 96636 7028 96692 7030
rect 96740 7082 96796 7084
rect 96740 7030 96742 7082
rect 96742 7030 96794 7082
rect 96794 7030 96796 7082
rect 96740 7028 96796 7030
rect 96844 7082 96900 7084
rect 96844 7030 96846 7082
rect 96846 7030 96898 7082
rect 96898 7030 96900 7082
rect 96844 7028 96900 7030
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 81276 6298 81332 6300
rect 81276 6246 81278 6298
rect 81278 6246 81330 6298
rect 81330 6246 81332 6298
rect 81276 6244 81332 6246
rect 81380 6298 81436 6300
rect 81380 6246 81382 6298
rect 81382 6246 81434 6298
rect 81434 6246 81436 6298
rect 81380 6244 81436 6246
rect 81484 6298 81540 6300
rect 81484 6246 81486 6298
rect 81486 6246 81538 6298
rect 81538 6246 81540 6298
rect 81484 6244 81540 6246
rect 111996 6298 112052 6300
rect 111996 6246 111998 6298
rect 111998 6246 112050 6298
rect 112050 6246 112052 6298
rect 111996 6244 112052 6246
rect 112100 6298 112156 6300
rect 112100 6246 112102 6298
rect 112102 6246 112154 6298
rect 112154 6246 112156 6298
rect 112100 6244 112156 6246
rect 112204 6298 112260 6300
rect 112204 6246 112206 6298
rect 112206 6246 112258 6298
rect 112258 6246 112260 6298
rect 112204 6244 112260 6246
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 96636 5514 96692 5516
rect 96636 5462 96638 5514
rect 96638 5462 96690 5514
rect 96690 5462 96692 5514
rect 96636 5460 96692 5462
rect 96740 5514 96796 5516
rect 96740 5462 96742 5514
rect 96742 5462 96794 5514
rect 96794 5462 96796 5514
rect 96740 5460 96796 5462
rect 96844 5514 96900 5516
rect 96844 5462 96846 5514
rect 96846 5462 96898 5514
rect 96898 5462 96900 5514
rect 96844 5460 96900 5462
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 81276 4730 81332 4732
rect 81276 4678 81278 4730
rect 81278 4678 81330 4730
rect 81330 4678 81332 4730
rect 81276 4676 81332 4678
rect 81380 4730 81436 4732
rect 81380 4678 81382 4730
rect 81382 4678 81434 4730
rect 81434 4678 81436 4730
rect 81380 4676 81436 4678
rect 81484 4730 81540 4732
rect 81484 4678 81486 4730
rect 81486 4678 81538 4730
rect 81538 4678 81540 4730
rect 81484 4676 81540 4678
rect 111996 4730 112052 4732
rect 111996 4678 111998 4730
rect 111998 4678 112050 4730
rect 112050 4678 112052 4730
rect 111996 4676 112052 4678
rect 112100 4730 112156 4732
rect 112100 4678 112102 4730
rect 112102 4678 112154 4730
rect 112154 4678 112156 4730
rect 112100 4676 112156 4678
rect 112204 4730 112260 4732
rect 112204 4678 112206 4730
rect 112206 4678 112258 4730
rect 112258 4678 112260 4730
rect 112204 4676 112260 4678
rect 20636 4172 20692 4228
rect 116508 4226 116564 4228
rect 116508 4174 116510 4226
rect 116510 4174 116562 4226
rect 116562 4174 116564 4226
rect 116508 4172 116564 4174
rect 116844 4172 116900 4228
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 96636 3946 96692 3948
rect 96636 3894 96638 3946
rect 96638 3894 96690 3946
rect 96690 3894 96692 3946
rect 96636 3892 96692 3894
rect 96740 3946 96796 3948
rect 96740 3894 96742 3946
rect 96742 3894 96794 3946
rect 96794 3894 96796 3946
rect 96740 3892 96796 3894
rect 96844 3946 96900 3948
rect 96844 3894 96846 3946
rect 96846 3894 96898 3946
rect 96898 3894 96900 3946
rect 96844 3892 96900 3894
rect 1820 2268 1876 2324
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 68572 3276 68628 3332
rect 69132 3330 69188 3332
rect 69132 3278 69134 3330
rect 69134 3278 69186 3330
rect 69186 3278 69188 3330
rect 69132 3276 69188 3278
rect 81276 3162 81332 3164
rect 81276 3110 81278 3162
rect 81278 3110 81330 3162
rect 81330 3110 81332 3162
rect 81276 3108 81332 3110
rect 81380 3162 81436 3164
rect 81380 3110 81382 3162
rect 81382 3110 81434 3162
rect 81434 3110 81436 3162
rect 81380 3108 81436 3110
rect 81484 3162 81540 3164
rect 81484 3110 81486 3162
rect 81486 3110 81538 3162
rect 81538 3110 81540 3162
rect 81484 3108 81540 3110
rect 106876 3276 106932 3332
rect 107660 3330 107716 3332
rect 107660 3278 107662 3330
rect 107662 3278 107714 3330
rect 107714 3278 107716 3330
rect 107660 3276 107716 3278
rect 111996 3162 112052 3164
rect 111996 3110 111998 3162
rect 111998 3110 112050 3162
rect 112050 3110 112052 3162
rect 111996 3108 112052 3110
rect 112100 3162 112156 3164
rect 112100 3110 112102 3162
rect 112102 3110 112154 3162
rect 112154 3110 112156 3162
rect 112100 3108 112156 3110
rect 112204 3162 112260 3164
rect 112204 3110 112206 3162
rect 112206 3110 112258 3162
rect 112258 3110 112260 3162
rect 112204 3108 112260 3110
rect 117740 3442 117796 3444
rect 117740 3390 117742 3442
rect 117742 3390 117794 3442
rect 117794 3390 117796 3442
rect 117740 3388 117796 3390
rect 118076 4060 118132 4116
rect 119644 3388 119700 3444
rect 117964 28 118020 84
<< metal3 >>
rect 200 135744 800 135856
rect 119200 135072 119800 135184
rect 200 134484 800 134512
rect 200 134428 2492 134484
rect 2548 134428 2558 134484
rect 200 134400 800 134428
rect 119200 133728 119800 133840
rect 200 133140 800 133168
rect 200 133084 1820 133140
rect 1876 133084 1886 133140
rect 200 133056 800 133084
rect 4466 132468 4476 132524
rect 4532 132468 4580 132524
rect 4636 132468 4684 132524
rect 4740 132468 4750 132524
rect 35186 132468 35196 132524
rect 35252 132468 35300 132524
rect 35356 132468 35404 132524
rect 35460 132468 35470 132524
rect 65906 132468 65916 132524
rect 65972 132468 66020 132524
rect 66076 132468 66124 132524
rect 66180 132468 66190 132524
rect 96626 132468 96636 132524
rect 96692 132468 96740 132524
rect 96796 132468 96844 132524
rect 96900 132468 96910 132524
rect 119200 132468 119800 132496
rect 117282 132412 117292 132468
rect 117348 132412 119800 132468
rect 119200 132384 119800 132412
rect 20178 132188 20188 132244
rect 20244 132188 22092 132244
rect 22148 132188 22158 132244
rect 59826 132076 59836 132132
rect 59892 132076 60844 132132
rect 60900 132076 60910 132132
rect 12786 131964 12796 132020
rect 12852 131964 13580 132020
rect 13636 131964 13646 132020
rect 71922 131964 71932 132020
rect 71988 131964 72380 132020
rect 72436 131964 72446 132020
rect 75282 131964 75292 132020
rect 75348 131964 76300 132020
rect 76356 131964 76366 132020
rect 95442 131964 95452 132020
rect 95508 131964 95900 132020
rect 95956 131964 95966 132020
rect 200 131712 800 131824
rect 19826 131684 19836 131740
rect 19892 131684 19940 131740
rect 19996 131684 20044 131740
rect 20100 131684 20110 131740
rect 50546 131684 50556 131740
rect 50612 131684 50660 131740
rect 50716 131684 50764 131740
rect 50820 131684 50830 131740
rect 81266 131684 81276 131740
rect 81332 131684 81380 131740
rect 81436 131684 81484 131740
rect 81540 131684 81550 131740
rect 111986 131684 111996 131740
rect 112052 131684 112100 131740
rect 112156 131684 112204 131740
rect 112260 131684 112270 131740
rect 119200 131040 119800 131152
rect 4466 130900 4476 130956
rect 4532 130900 4580 130956
rect 4636 130900 4684 130956
rect 4740 130900 4750 130956
rect 35186 130900 35196 130956
rect 35252 130900 35300 130956
rect 35356 130900 35404 130956
rect 35460 130900 35470 130956
rect 65906 130900 65916 130956
rect 65972 130900 66020 130956
rect 66076 130900 66124 130956
rect 66180 130900 66190 130956
rect 96626 130900 96636 130956
rect 96692 130900 96740 130956
rect 96796 130900 96844 130956
rect 96900 130900 96910 130956
rect 200 130452 800 130480
rect 200 130396 1820 130452
rect 1876 130396 1886 130452
rect 200 130368 800 130396
rect 19826 130116 19836 130172
rect 19892 130116 19940 130172
rect 19996 130116 20044 130172
rect 20100 130116 20110 130172
rect 50546 130116 50556 130172
rect 50612 130116 50660 130172
rect 50716 130116 50764 130172
rect 50820 130116 50830 130172
rect 81266 130116 81276 130172
rect 81332 130116 81380 130172
rect 81436 130116 81484 130172
rect 81540 130116 81550 130172
rect 111986 130116 111996 130172
rect 112052 130116 112100 130172
rect 112156 130116 112204 130172
rect 112260 130116 112270 130172
rect 119200 129696 119800 129808
rect 4466 129332 4476 129388
rect 4532 129332 4580 129388
rect 4636 129332 4684 129388
rect 4740 129332 4750 129388
rect 35186 129332 35196 129388
rect 35252 129332 35300 129388
rect 35356 129332 35404 129388
rect 35460 129332 35470 129388
rect 65906 129332 65916 129388
rect 65972 129332 66020 129388
rect 66076 129332 66124 129388
rect 66180 129332 66190 129388
rect 96626 129332 96636 129388
rect 96692 129332 96740 129388
rect 96796 129332 96844 129388
rect 96900 129332 96910 129388
rect 200 129024 800 129136
rect 19826 128548 19836 128604
rect 19892 128548 19940 128604
rect 19996 128548 20044 128604
rect 20100 128548 20110 128604
rect 50546 128548 50556 128604
rect 50612 128548 50660 128604
rect 50716 128548 50764 128604
rect 50820 128548 50830 128604
rect 81266 128548 81276 128604
rect 81332 128548 81380 128604
rect 81436 128548 81484 128604
rect 81540 128548 81550 128604
rect 111986 128548 111996 128604
rect 112052 128548 112100 128604
rect 112156 128548 112204 128604
rect 112260 128548 112270 128604
rect 119200 128352 119800 128464
rect 200 127764 800 127792
rect 4466 127764 4476 127820
rect 4532 127764 4580 127820
rect 4636 127764 4684 127820
rect 4740 127764 4750 127820
rect 35186 127764 35196 127820
rect 35252 127764 35300 127820
rect 35356 127764 35404 127820
rect 35460 127764 35470 127820
rect 65906 127764 65916 127820
rect 65972 127764 66020 127820
rect 66076 127764 66124 127820
rect 66180 127764 66190 127820
rect 96626 127764 96636 127820
rect 96692 127764 96740 127820
rect 96796 127764 96844 127820
rect 96900 127764 96910 127820
rect 200 127708 1820 127764
rect 1876 127708 1886 127764
rect 200 127680 800 127708
rect 119200 127680 119800 127792
rect 200 127092 800 127120
rect 200 127036 1820 127092
rect 1876 127036 1886 127092
rect 200 127008 800 127036
rect 19826 126980 19836 127036
rect 19892 126980 19940 127036
rect 19996 126980 20044 127036
rect 20100 126980 20110 127036
rect 50546 126980 50556 127036
rect 50612 126980 50660 127036
rect 50716 126980 50764 127036
rect 50820 126980 50830 127036
rect 81266 126980 81276 127036
rect 81332 126980 81380 127036
rect 81436 126980 81484 127036
rect 81540 126980 81550 127036
rect 111986 126980 111996 127036
rect 112052 126980 112100 127036
rect 112156 126980 112204 127036
rect 112260 126980 112270 127036
rect 119200 126420 119800 126448
rect 118066 126364 118076 126420
rect 118132 126364 119800 126420
rect 119200 126336 119800 126364
rect 4466 126196 4476 126252
rect 4532 126196 4580 126252
rect 4636 126196 4684 126252
rect 4740 126196 4750 126252
rect 35186 126196 35196 126252
rect 35252 126196 35300 126252
rect 35356 126196 35404 126252
rect 35460 126196 35470 126252
rect 65906 126196 65916 126252
rect 65972 126196 66020 126252
rect 66076 126196 66124 126252
rect 66180 126196 66190 126252
rect 96626 126196 96636 126252
rect 96692 126196 96740 126252
rect 96796 126196 96844 126252
rect 96900 126196 96910 126252
rect 200 125664 800 125776
rect 19826 125412 19836 125468
rect 19892 125412 19940 125468
rect 19996 125412 20044 125468
rect 20100 125412 20110 125468
rect 50546 125412 50556 125468
rect 50612 125412 50660 125468
rect 50716 125412 50764 125468
rect 50820 125412 50830 125468
rect 81266 125412 81276 125468
rect 81332 125412 81380 125468
rect 81436 125412 81484 125468
rect 81540 125412 81550 125468
rect 111986 125412 111996 125468
rect 112052 125412 112100 125468
rect 112156 125412 112204 125468
rect 112260 125412 112270 125468
rect 119200 124992 119800 125104
rect 4466 124628 4476 124684
rect 4532 124628 4580 124684
rect 4636 124628 4684 124684
rect 4740 124628 4750 124684
rect 35186 124628 35196 124684
rect 35252 124628 35300 124684
rect 35356 124628 35404 124684
rect 35460 124628 35470 124684
rect 65906 124628 65916 124684
rect 65972 124628 66020 124684
rect 66076 124628 66124 124684
rect 66180 124628 66190 124684
rect 96626 124628 96636 124684
rect 96692 124628 96740 124684
rect 96796 124628 96844 124684
rect 96900 124628 96910 124684
rect 200 124404 800 124432
rect 200 124348 1820 124404
rect 1876 124348 1886 124404
rect 200 124320 800 124348
rect 19826 123844 19836 123900
rect 19892 123844 19940 123900
rect 19996 123844 20044 123900
rect 20100 123844 20110 123900
rect 50546 123844 50556 123900
rect 50612 123844 50660 123900
rect 50716 123844 50764 123900
rect 50820 123844 50830 123900
rect 81266 123844 81276 123900
rect 81332 123844 81380 123900
rect 81436 123844 81484 123900
rect 81540 123844 81550 123900
rect 111986 123844 111996 123900
rect 112052 123844 112100 123900
rect 112156 123844 112204 123900
rect 112260 123844 112270 123900
rect 119200 123732 119800 123760
rect 118066 123676 118076 123732
rect 118132 123676 119800 123732
rect 119200 123648 119800 123676
rect 200 123060 800 123088
rect 4466 123060 4476 123116
rect 4532 123060 4580 123116
rect 4636 123060 4684 123116
rect 4740 123060 4750 123116
rect 35186 123060 35196 123116
rect 35252 123060 35300 123116
rect 35356 123060 35404 123116
rect 35460 123060 35470 123116
rect 65906 123060 65916 123116
rect 65972 123060 66020 123116
rect 66076 123060 66124 123116
rect 66180 123060 66190 123116
rect 96626 123060 96636 123116
rect 96692 123060 96740 123116
rect 96796 123060 96844 123116
rect 96900 123060 96910 123116
rect 200 123004 1820 123060
rect 1876 123004 1886 123060
rect 200 122976 800 123004
rect 19826 122276 19836 122332
rect 19892 122276 19940 122332
rect 19996 122276 20044 122332
rect 20100 122276 20110 122332
rect 50546 122276 50556 122332
rect 50612 122276 50660 122332
rect 50716 122276 50764 122332
rect 50820 122276 50830 122332
rect 81266 122276 81276 122332
rect 81332 122276 81380 122332
rect 81436 122276 81484 122332
rect 81540 122276 81550 122332
rect 111986 122276 111996 122332
rect 112052 122276 112100 122332
rect 112156 122276 112204 122332
rect 112260 122276 112270 122332
rect 119200 122304 119800 122416
rect 200 121716 800 121744
rect 200 121660 1820 121716
rect 1876 121660 1886 121716
rect 200 121632 800 121660
rect 4466 121492 4476 121548
rect 4532 121492 4580 121548
rect 4636 121492 4684 121548
rect 4740 121492 4750 121548
rect 35186 121492 35196 121548
rect 35252 121492 35300 121548
rect 35356 121492 35404 121548
rect 35460 121492 35470 121548
rect 65906 121492 65916 121548
rect 65972 121492 66020 121548
rect 66076 121492 66124 121548
rect 66180 121492 66190 121548
rect 96626 121492 96636 121548
rect 96692 121492 96740 121548
rect 96796 121492 96844 121548
rect 96900 121492 96910 121548
rect 119200 120960 119800 121072
rect 19826 120708 19836 120764
rect 19892 120708 19940 120764
rect 19996 120708 20044 120764
rect 20100 120708 20110 120764
rect 50546 120708 50556 120764
rect 50612 120708 50660 120764
rect 50716 120708 50764 120764
rect 50820 120708 50830 120764
rect 81266 120708 81276 120764
rect 81332 120708 81380 120764
rect 81436 120708 81484 120764
rect 81540 120708 81550 120764
rect 111986 120708 111996 120764
rect 112052 120708 112100 120764
rect 112156 120708 112204 120764
rect 112260 120708 112270 120764
rect 200 120288 800 120400
rect 119200 120288 119800 120400
rect 4466 119924 4476 119980
rect 4532 119924 4580 119980
rect 4636 119924 4684 119980
rect 4740 119924 4750 119980
rect 35186 119924 35196 119980
rect 35252 119924 35300 119980
rect 35356 119924 35404 119980
rect 35460 119924 35470 119980
rect 65906 119924 65916 119980
rect 65972 119924 66020 119980
rect 66076 119924 66124 119980
rect 66180 119924 66190 119980
rect 96626 119924 96636 119980
rect 96692 119924 96740 119980
rect 96796 119924 96844 119980
rect 96900 119924 96910 119980
rect 200 119616 800 119728
rect 19826 119140 19836 119196
rect 19892 119140 19940 119196
rect 19996 119140 20044 119196
rect 20100 119140 20110 119196
rect 50546 119140 50556 119196
rect 50612 119140 50660 119196
rect 50716 119140 50764 119196
rect 50820 119140 50830 119196
rect 81266 119140 81276 119196
rect 81332 119140 81380 119196
rect 81436 119140 81484 119196
rect 81540 119140 81550 119196
rect 111986 119140 111996 119196
rect 112052 119140 112100 119196
rect 112156 119140 112204 119196
rect 112260 119140 112270 119196
rect 119200 118944 119800 119056
rect 200 118272 800 118384
rect 4466 118356 4476 118412
rect 4532 118356 4580 118412
rect 4636 118356 4684 118412
rect 4740 118356 4750 118412
rect 35186 118356 35196 118412
rect 35252 118356 35300 118412
rect 35356 118356 35404 118412
rect 35460 118356 35470 118412
rect 65906 118356 65916 118412
rect 65972 118356 66020 118412
rect 66076 118356 66124 118412
rect 66180 118356 66190 118412
rect 96626 118356 96636 118412
rect 96692 118356 96740 118412
rect 96796 118356 96844 118412
rect 96900 118356 96910 118412
rect 19826 117572 19836 117628
rect 19892 117572 19940 117628
rect 19996 117572 20044 117628
rect 20100 117572 20110 117628
rect 50546 117572 50556 117628
rect 50612 117572 50660 117628
rect 50716 117572 50764 117628
rect 50820 117572 50830 117628
rect 81266 117572 81276 117628
rect 81332 117572 81380 117628
rect 81436 117572 81484 117628
rect 81540 117572 81550 117628
rect 111986 117572 111996 117628
rect 112052 117572 112100 117628
rect 112156 117572 112204 117628
rect 112260 117572 112270 117628
rect 119200 117600 119800 117712
rect 200 117012 800 117040
rect 200 116956 1820 117012
rect 1876 116956 1886 117012
rect 200 116928 800 116956
rect 4466 116788 4476 116844
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4740 116788 4750 116844
rect 35186 116788 35196 116844
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35460 116788 35470 116844
rect 65906 116788 65916 116844
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 66180 116788 66190 116844
rect 96626 116788 96636 116844
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96900 116788 96910 116844
rect 119200 116340 119800 116368
rect 118066 116284 118076 116340
rect 118132 116284 119800 116340
rect 119200 116256 119800 116284
rect 19826 116004 19836 116060
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 20100 116004 20110 116060
rect 50546 116004 50556 116060
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50820 116004 50830 116060
rect 81266 116004 81276 116060
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81540 116004 81550 116060
rect 111986 116004 111996 116060
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 112260 116004 112270 116060
rect 200 115584 800 115696
rect 4466 115220 4476 115276
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4740 115220 4750 115276
rect 35186 115220 35196 115276
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35460 115220 35470 115276
rect 65906 115220 65916 115276
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 66180 115220 66190 115276
rect 96626 115220 96636 115276
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96900 115220 96910 115276
rect 119200 114996 119800 115024
rect 118066 114940 118076 114996
rect 118132 114940 119800 114996
rect 119200 114912 119800 114940
rect 19826 114436 19836 114492
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 20100 114436 20110 114492
rect 50546 114436 50556 114492
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50820 114436 50830 114492
rect 81266 114436 81276 114492
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81540 114436 81550 114492
rect 111986 114436 111996 114492
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 112260 114436 112270 114492
rect 200 114240 800 114352
rect 4466 113652 4476 113708
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4740 113652 4750 113708
rect 35186 113652 35196 113708
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35460 113652 35470 113708
rect 65906 113652 65916 113708
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 66180 113652 66190 113708
rect 96626 113652 96636 113708
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96900 113652 96910 113708
rect 119200 113652 119800 113680
rect 117618 113596 117628 113652
rect 117684 113596 119800 113652
rect 119200 113568 119800 113596
rect 200 112896 800 113008
rect 19826 112868 19836 112924
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 20100 112868 20110 112924
rect 50546 112868 50556 112924
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50820 112868 50830 112924
rect 81266 112868 81276 112924
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81540 112868 81550 112924
rect 111986 112868 111996 112924
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 112260 112868 112270 112924
rect 119200 112896 119800 113008
rect 200 112224 800 112336
rect 4466 112084 4476 112140
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4740 112084 4750 112140
rect 35186 112084 35196 112140
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35460 112084 35470 112140
rect 65906 112084 65916 112140
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 66180 112084 66190 112140
rect 96626 112084 96636 112140
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96900 112084 96910 112140
rect 119200 111636 119800 111664
rect 118066 111580 118076 111636
rect 118132 111580 119800 111636
rect 119200 111552 119800 111580
rect 19826 111300 19836 111356
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 20100 111300 20110 111356
rect 50546 111300 50556 111356
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50820 111300 50830 111356
rect 81266 111300 81276 111356
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81540 111300 81550 111356
rect 111986 111300 111996 111356
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 112260 111300 112270 111356
rect 200 110964 800 110992
rect 200 110908 1820 110964
rect 1876 110908 1886 110964
rect 200 110880 800 110908
rect 4466 110516 4476 110572
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4740 110516 4750 110572
rect 35186 110516 35196 110572
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35460 110516 35470 110572
rect 65906 110516 65916 110572
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 66180 110516 66190 110572
rect 96626 110516 96636 110572
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96900 110516 96910 110572
rect 119200 110292 119800 110320
rect 118066 110236 118076 110292
rect 118132 110236 119800 110292
rect 119200 110208 119800 110236
rect 19826 109732 19836 109788
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 20100 109732 20110 109788
rect 50546 109732 50556 109788
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50820 109732 50830 109788
rect 81266 109732 81276 109788
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81540 109732 81550 109788
rect 111986 109732 111996 109788
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 112260 109732 112270 109788
rect 200 109620 800 109648
rect 200 109564 1820 109620
rect 1876 109564 1886 109620
rect 200 109536 800 109564
rect 4466 108948 4476 109004
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4740 108948 4750 109004
rect 35186 108948 35196 109004
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35460 108948 35470 109004
rect 65906 108948 65916 109004
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 66180 108948 66190 109004
rect 96626 108948 96636 109004
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96900 108948 96910 109004
rect 119200 108864 119800 108976
rect 200 108192 800 108304
rect 19826 108164 19836 108220
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 20100 108164 20110 108220
rect 50546 108164 50556 108220
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50820 108164 50830 108220
rect 81266 108164 81276 108220
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81540 108164 81550 108220
rect 111986 108164 111996 108220
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 112260 108164 112270 108220
rect 119200 107604 119800 107632
rect 118066 107548 118076 107604
rect 118132 107548 119800 107604
rect 119200 107520 119800 107548
rect 4466 107380 4476 107436
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4740 107380 4750 107436
rect 35186 107380 35196 107436
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35460 107380 35470 107436
rect 65906 107380 65916 107436
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 66180 107380 66190 107436
rect 96626 107380 96636 107436
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96900 107380 96910 107436
rect 200 106848 800 106960
rect 19826 106596 19836 106652
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 20100 106596 20110 106652
rect 50546 106596 50556 106652
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50820 106596 50830 106652
rect 81266 106596 81276 106652
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81540 106596 81550 106652
rect 111986 106596 111996 106652
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 112260 106596 112270 106652
rect 119200 106260 119800 106288
rect 118066 106204 118076 106260
rect 118132 106204 119800 106260
rect 119200 106176 119800 106204
rect 4466 105812 4476 105868
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4740 105812 4750 105868
rect 35186 105812 35196 105868
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35460 105812 35470 105868
rect 65906 105812 65916 105868
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 66180 105812 66190 105868
rect 96626 105812 96636 105868
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96900 105812 96910 105868
rect 200 105504 800 105616
rect 119200 105504 119800 105616
rect 19826 105028 19836 105084
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 20100 105028 20110 105084
rect 50546 105028 50556 105084
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50820 105028 50830 105084
rect 81266 105028 81276 105084
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81540 105028 81550 105084
rect 111986 105028 111996 105084
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 112260 105028 112270 105084
rect 200 104916 800 104944
rect 200 104860 1820 104916
rect 1876 104860 1886 104916
rect 200 104832 800 104860
rect 4466 104244 4476 104300
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4740 104244 4750 104300
rect 35186 104244 35196 104300
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35460 104244 35470 104300
rect 65906 104244 65916 104300
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 66180 104244 66190 104300
rect 96626 104244 96636 104300
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96900 104244 96910 104300
rect 119200 104160 119800 104272
rect 200 103488 800 103600
rect 19826 103460 19836 103516
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 20100 103460 20110 103516
rect 50546 103460 50556 103516
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50820 103460 50830 103516
rect 81266 103460 81276 103516
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81540 103460 81550 103516
rect 111986 103460 111996 103516
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 112260 103460 112270 103516
rect 119200 102900 119800 102928
rect 118066 102844 118076 102900
rect 118132 102844 119800 102900
rect 119200 102816 119800 102844
rect 4466 102676 4476 102732
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4740 102676 4750 102732
rect 35186 102676 35196 102732
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35460 102676 35470 102732
rect 65906 102676 65916 102732
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 66180 102676 66190 102732
rect 96626 102676 96636 102732
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96900 102676 96910 102732
rect 200 102144 800 102256
rect 19826 101892 19836 101948
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 20100 101892 20110 101948
rect 50546 101892 50556 101948
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50820 101892 50830 101948
rect 81266 101892 81276 101948
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81540 101892 81550 101948
rect 111986 101892 111996 101948
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 112260 101892 112270 101948
rect 119200 101472 119800 101584
rect 4466 101108 4476 101164
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4740 101108 4750 101164
rect 35186 101108 35196 101164
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35460 101108 35470 101164
rect 65906 101108 65916 101164
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 66180 101108 66190 101164
rect 96626 101108 96636 101164
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96900 101108 96910 101164
rect 200 100884 800 100912
rect 200 100828 1820 100884
rect 1876 100828 1886 100884
rect 200 100800 800 100828
rect 19826 100324 19836 100380
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 20100 100324 20110 100380
rect 50546 100324 50556 100380
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50820 100324 50830 100380
rect 81266 100324 81276 100380
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81540 100324 81550 100380
rect 111986 100324 111996 100380
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 112260 100324 112270 100380
rect 119200 100128 119800 100240
rect 200 99456 800 99568
rect 4466 99540 4476 99596
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4740 99540 4750 99596
rect 35186 99540 35196 99596
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35460 99540 35470 99596
rect 65906 99540 65916 99596
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 66180 99540 66190 99596
rect 96626 99540 96636 99596
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96900 99540 96910 99596
rect 19826 98756 19836 98812
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 20100 98756 20110 98812
rect 50546 98756 50556 98812
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50820 98756 50830 98812
rect 81266 98756 81276 98812
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81540 98756 81550 98812
rect 111986 98756 111996 98812
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 112260 98756 112270 98812
rect 119200 98784 119800 98896
rect 200 98112 800 98224
rect 119200 98196 119800 98224
rect 118066 98140 118076 98196
rect 118132 98140 119800 98196
rect 119200 98112 119800 98140
rect 4466 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4750 98028
rect 35186 97972 35196 98028
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35460 97972 35470 98028
rect 65906 97972 65916 98028
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 66180 97972 66190 98028
rect 96626 97972 96636 98028
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96900 97972 96910 98028
rect 200 97440 800 97552
rect 19826 97188 19836 97244
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 20100 97188 20110 97244
rect 50546 97188 50556 97244
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50820 97188 50830 97244
rect 81266 97188 81276 97244
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81540 97188 81550 97244
rect 111986 97188 111996 97244
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 112260 97188 112270 97244
rect 119200 96852 119800 96880
rect 118066 96796 118076 96852
rect 118132 96796 119800 96852
rect 119200 96768 119800 96796
rect 4466 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4750 96460
rect 35186 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35470 96460
rect 65906 96404 65916 96460
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 66180 96404 66190 96460
rect 96626 96404 96636 96460
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96900 96404 96910 96460
rect 200 96180 800 96208
rect 200 96124 1820 96180
rect 1876 96124 1886 96180
rect 200 96096 800 96124
rect 19826 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20110 95676
rect 50546 95620 50556 95676
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50820 95620 50830 95676
rect 81266 95620 81276 95676
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81540 95620 81550 95676
rect 111986 95620 111996 95676
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 112260 95620 112270 95676
rect 119200 95508 119800 95536
rect 118066 95452 118076 95508
rect 118132 95452 119800 95508
rect 119200 95424 119800 95452
rect 200 94836 800 94864
rect 4466 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4750 94892
rect 35186 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35470 94892
rect 65906 94836 65916 94892
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 66180 94836 66190 94892
rect 96626 94836 96636 94892
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96900 94836 96910 94892
rect 200 94780 1820 94836
rect 1876 94780 1886 94836
rect 200 94752 800 94780
rect 19826 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20110 94108
rect 50546 94052 50556 94108
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50820 94052 50830 94108
rect 81266 94052 81276 94108
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81540 94052 81550 94108
rect 111986 94052 111996 94108
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 112260 94052 112270 94108
rect 119200 94080 119800 94192
rect 200 93408 800 93520
rect 4466 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4750 93324
rect 35186 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35470 93324
rect 65906 93268 65916 93324
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 66180 93268 66190 93324
rect 96626 93268 96636 93324
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96900 93268 96910 93324
rect 119200 92736 119800 92848
rect 19826 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20110 92540
rect 50546 92484 50556 92540
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50820 92484 50830 92540
rect 81266 92484 81276 92540
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81540 92484 81550 92540
rect 111986 92484 111996 92540
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 112260 92484 112270 92540
rect 200 92148 800 92176
rect 200 92092 1820 92148
rect 1876 92092 1886 92148
rect 200 92064 800 92092
rect 4466 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4750 91756
rect 35186 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35470 91756
rect 65906 91700 65916 91756
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 66180 91700 66190 91756
rect 96626 91700 96636 91756
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96900 91700 96910 91756
rect 119200 91392 119800 91504
rect 19826 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20110 90972
rect 50546 90916 50556 90972
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50820 90916 50830 90972
rect 81266 90916 81276 90972
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81540 90916 81550 90972
rect 111986 90916 111996 90972
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 112260 90916 112270 90972
rect 200 90804 800 90832
rect 119200 90804 119800 90832
rect 200 90748 1820 90804
rect 1876 90748 1886 90804
rect 118066 90748 118076 90804
rect 118132 90748 119800 90804
rect 200 90720 800 90748
rect 119200 90720 119800 90748
rect 200 90132 800 90160
rect 4466 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4750 90188
rect 35186 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35470 90188
rect 65906 90132 65916 90188
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 66180 90132 66190 90188
rect 96626 90132 96636 90188
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96900 90132 96910 90188
rect 200 90076 1820 90132
rect 1876 90076 1886 90132
rect 200 90048 800 90076
rect 19826 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20110 89404
rect 50546 89348 50556 89404
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50820 89348 50830 89404
rect 81266 89348 81276 89404
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81540 89348 81550 89404
rect 111986 89348 111996 89404
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 112260 89348 112270 89404
rect 119200 89376 119800 89488
rect 200 88704 800 88816
rect 4466 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4750 88620
rect 35186 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35470 88620
rect 65906 88564 65916 88620
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 66180 88564 66190 88620
rect 96626 88564 96636 88620
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96900 88564 96910 88620
rect 119200 88116 119800 88144
rect 118066 88060 118076 88116
rect 118132 88060 119800 88116
rect 119200 88032 119800 88060
rect 19826 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20110 87836
rect 50546 87780 50556 87836
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50820 87780 50830 87836
rect 81266 87780 81276 87836
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81540 87780 81550 87836
rect 111986 87780 111996 87836
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 112260 87780 112270 87836
rect 200 87360 800 87472
rect 4466 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4750 87052
rect 35186 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35470 87052
rect 65906 86996 65916 87052
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 66180 86996 66190 87052
rect 96626 86996 96636 87052
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96900 86996 96910 87052
rect 119200 86688 119800 86800
rect 19826 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20110 86268
rect 50546 86212 50556 86268
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50820 86212 50830 86268
rect 81266 86212 81276 86268
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81540 86212 81550 86268
rect 111986 86212 111996 86268
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 112260 86212 112270 86268
rect 200 86016 800 86128
rect 4466 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4750 85484
rect 35186 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35470 85484
rect 65906 85428 65916 85484
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 66180 85428 66190 85484
rect 96626 85428 96636 85484
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96900 85428 96910 85484
rect 119200 85344 119800 85456
rect 2818 84812 2828 84868
rect 2884 84812 3500 84868
rect 3556 84812 3566 84868
rect 200 84756 800 84784
rect 200 84700 2156 84756
rect 2212 84700 2222 84756
rect 200 84672 800 84700
rect 19826 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20110 84700
rect 50546 84644 50556 84700
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50820 84644 50830 84700
rect 81266 84644 81276 84700
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81540 84644 81550 84700
rect 111986 84644 111996 84700
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 112260 84644 112270 84700
rect 119200 84084 119800 84112
rect 118066 84028 118076 84084
rect 118132 84028 119800 84084
rect 119200 84000 119800 84028
rect 4466 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4750 83916
rect 35186 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35470 83916
rect 65906 83860 65916 83916
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 66180 83860 66190 83916
rect 96626 83860 96636 83916
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96900 83860 96910 83916
rect 200 83412 800 83440
rect 200 83356 2492 83412
rect 2548 83356 2558 83412
rect 200 83328 800 83356
rect 119200 83328 119800 83440
rect 19826 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20110 83132
rect 50546 83076 50556 83132
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50820 83076 50830 83132
rect 81266 83076 81276 83132
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81540 83076 81550 83132
rect 111986 83076 111996 83132
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 112260 83076 112270 83132
rect 200 82740 800 82768
rect 200 82684 1820 82740
rect 1876 82684 1886 82740
rect 200 82656 800 82684
rect 4466 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4750 82348
rect 35186 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35470 82348
rect 65906 82292 65916 82348
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 66180 82292 66190 82348
rect 96626 82292 96636 82348
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96900 82292 96910 82348
rect 119200 82068 119800 82096
rect 118066 82012 118076 82068
rect 118132 82012 119800 82068
rect 119200 81984 119800 82012
rect 19826 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20110 81564
rect 50546 81508 50556 81564
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50820 81508 50830 81564
rect 81266 81508 81276 81564
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81540 81508 81550 81564
rect 111986 81508 111996 81564
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 112260 81508 112270 81564
rect 200 81312 800 81424
rect 4466 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4750 80780
rect 35186 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35470 80780
rect 65906 80724 65916 80780
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 66180 80724 66190 80780
rect 96626 80724 96636 80780
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96900 80724 96910 80780
rect 119200 80640 119800 80752
rect 200 79968 800 80080
rect 19826 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20110 79996
rect 50546 79940 50556 79996
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50820 79940 50830 79996
rect 81266 79940 81276 79996
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81540 79940 81550 79996
rect 111986 79940 111996 79996
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 112260 79940 112270 79996
rect 119200 79380 119800 79408
rect 118066 79324 118076 79380
rect 118132 79324 119800 79380
rect 119200 79296 119800 79324
rect 4466 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4750 79212
rect 35186 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35470 79212
rect 65906 79156 65916 79212
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 66180 79156 66190 79212
rect 96626 79156 96636 79212
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96900 79156 96910 79212
rect 200 78624 800 78736
rect 19826 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20110 78428
rect 50546 78372 50556 78428
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50820 78372 50830 78428
rect 81266 78372 81276 78428
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81540 78372 81550 78428
rect 111986 78372 111996 78428
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 112260 78372 112270 78428
rect 119200 77952 119800 78064
rect 4466 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4750 77644
rect 35186 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35470 77644
rect 65906 77588 65916 77644
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 66180 77588 66190 77644
rect 96626 77588 96636 77644
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96900 77588 96910 77644
rect 200 77364 800 77392
rect 200 77308 1820 77364
rect 1876 77308 1886 77364
rect 200 77280 800 77308
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 81266 76804 81276 76860
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81540 76804 81550 76860
rect 111986 76804 111996 76860
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 112260 76804 112270 76860
rect 119200 76692 119800 76720
rect 118066 76636 118076 76692
rect 118132 76636 119800 76692
rect 119200 76608 119800 76636
rect 200 75936 800 76048
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 96626 76020 96636 76076
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96900 76020 96910 76076
rect 119200 75936 119800 76048
rect 200 75264 800 75376
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 81266 75236 81276 75292
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81540 75236 81550 75292
rect 111986 75236 111996 75292
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 112260 75236 112270 75292
rect 119200 74592 119800 74704
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 96626 74452 96636 74508
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96900 74452 96910 74508
rect 200 73920 800 74032
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 81266 73668 81276 73724
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81540 73668 81550 73724
rect 111986 73668 111996 73724
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 112260 73668 112270 73724
rect 119200 73332 119800 73360
rect 118066 73276 118076 73332
rect 118132 73276 119800 73332
rect 119200 73248 119800 73276
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 96626 72884 96636 72940
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96900 72884 96910 72940
rect 200 72660 800 72688
rect 200 72604 1820 72660
rect 1876 72604 1886 72660
rect 200 72576 800 72604
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 81266 72100 81276 72156
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81540 72100 81550 72156
rect 111986 72100 111996 72156
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 112260 72100 112270 72156
rect 119200 71904 119800 72016
rect 200 71232 800 71344
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 96626 71316 96636 71372
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96900 71316 96910 71372
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 81266 70532 81276 70588
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81540 70532 81550 70588
rect 111986 70532 111996 70588
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 112260 70532 112270 70588
rect 119200 70560 119800 70672
rect 200 69888 800 70000
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 96626 69748 96636 69804
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96900 69748 96910 69804
rect 119200 69300 119800 69328
rect 118066 69244 118076 69300
rect 118132 69244 119800 69300
rect 119200 69216 119800 69244
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 81266 68964 81276 69020
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81540 68964 81550 69020
rect 111986 68964 111996 69020
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 112260 68964 112270 69020
rect 2594 68796 2604 68852
rect 2660 68796 3164 68852
rect 3220 68796 3230 68852
rect 20066 68796 20076 68852
rect 20132 68796 21420 68852
rect 21476 68796 21486 68852
rect 200 68544 800 68656
rect 19954 68460 19964 68516
rect 20020 68460 20636 68516
rect 20692 68460 20702 68516
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 96626 68180 96636 68236
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96900 68180 96910 68236
rect 200 67872 800 67984
rect 119200 67956 119800 67984
rect 59602 67900 59612 67956
rect 59668 67900 60060 67956
rect 60116 67900 60620 67956
rect 60676 67900 60686 67956
rect 118066 67900 118076 67956
rect 118132 67900 119800 67956
rect 119200 67872 119800 67900
rect 2706 67564 2716 67620
rect 2772 67564 3500 67620
rect 3556 67564 5068 67620
rect 5124 67564 5134 67620
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 81266 67396 81276 67452
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81540 67396 81550 67452
rect 111986 67396 111996 67452
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 112260 67396 112270 67452
rect 119200 67284 119800 67312
rect 118066 67228 118076 67284
rect 118132 67228 119800 67284
rect 119200 67200 119800 67228
rect 1922 67116 1932 67172
rect 1988 67116 6300 67172
rect 6356 67116 6366 67172
rect 3714 67004 3724 67060
rect 3780 67004 4620 67060
rect 4676 67004 4686 67060
rect 5842 66780 5852 66836
rect 5908 66780 20636 66836
rect 20692 66780 20702 66836
rect 200 66612 800 66640
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 96626 66612 96636 66668
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96900 66612 96910 66668
rect 200 66556 1820 66612
rect 1876 66556 1886 66612
rect 200 66528 800 66556
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 81266 65828 81276 65884
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81540 65828 81550 65884
rect 111986 65828 111996 65884
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 112260 65828 112270 65884
rect 119200 65856 119800 65968
rect 200 65184 800 65296
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 96626 65044 96636 65100
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96900 65044 96910 65100
rect 119200 64512 119800 64624
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 81266 64260 81276 64316
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81540 64260 81550 64316
rect 111986 64260 111996 64316
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 112260 64260 112270 64316
rect 200 63924 800 63952
rect 200 63868 1820 63924
rect 1876 63868 1886 63924
rect 200 63840 800 63868
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 96626 63476 96636 63532
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96900 63476 96910 63532
rect 119200 63168 119800 63280
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 81266 62692 81276 62748
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81540 62692 81550 62748
rect 111986 62692 111996 62748
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 112260 62692 112270 62748
rect 200 62496 800 62608
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 96626 61908 96636 61964
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96900 61908 96910 61964
rect 119200 61824 119800 61936
rect 200 61236 800 61264
rect 200 61180 1820 61236
rect 1876 61180 1886 61236
rect 200 61152 800 61180
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 81266 61124 81276 61180
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81540 61124 81550 61180
rect 111986 61124 111996 61180
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 112260 61124 112270 61180
rect 119200 60564 119800 60592
rect 118066 60508 118076 60564
rect 118132 60508 119800 60564
rect 119200 60480 119800 60508
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 96626 60340 96636 60396
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96900 60340 96910 60396
rect 200 59808 800 59920
rect 119200 59892 119800 59920
rect 118066 59836 118076 59892
rect 118132 59836 119800 59892
rect 119200 59808 119800 59836
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 81266 59556 81276 59612
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81540 59556 81550 59612
rect 111986 59556 111996 59612
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 112260 59556 112270 59612
rect 200 59136 800 59248
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 96626 58772 96636 58828
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96900 58772 96910 58828
rect 119200 58548 119800 58576
rect 118066 58492 118076 58548
rect 118132 58492 119800 58548
rect 119200 58464 119800 58492
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 81266 57988 81276 58044
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81540 57988 81550 58044
rect 111986 57988 111996 58044
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 112260 57988 112270 58044
rect 200 57876 800 57904
rect 200 57820 1820 57876
rect 1876 57820 1886 57876
rect 200 57792 800 57820
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 96626 57204 96636 57260
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96900 57204 96910 57260
rect 119200 57204 119800 57232
rect 118066 57148 118076 57204
rect 118132 57148 119800 57204
rect 119200 57120 119800 57148
rect 200 56448 800 56560
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 81266 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81550 56476
rect 111986 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112270 56476
rect 119200 55776 119800 55888
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 96626 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96910 55692
rect 200 55104 800 55216
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 81266 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81550 54908
rect 111986 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112270 54908
rect 119200 54432 119800 54544
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 96626 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96910 54124
rect 200 53760 800 53872
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 81266 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81550 53340
rect 111986 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112270 53340
rect 118066 53228 118076 53284
rect 118132 53228 118142 53284
rect 118076 53172 118132 53228
rect 119200 53172 119800 53200
rect 118076 53116 119800 53172
rect 119200 53088 119800 53116
rect 200 52500 800 52528
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 96626 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96910 52556
rect 119200 52500 119800 52528
rect 200 52444 1820 52500
rect 1876 52444 1886 52500
rect 118066 52444 118076 52500
rect 118132 52444 119800 52500
rect 200 52416 800 52444
rect 119200 52416 119800 52444
rect 200 51744 800 51856
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 81266 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81550 51772
rect 111986 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112270 51772
rect 119200 51072 119800 51184
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 96626 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96910 50988
rect 200 50400 800 50512
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 81266 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81550 50204
rect 111986 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112270 50204
rect 119200 49728 119800 49840
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 96626 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96910 49420
rect 200 49140 800 49168
rect 200 49084 1820 49140
rect 1876 49084 1886 49140
rect 200 49056 800 49084
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 81266 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81550 48636
rect 111986 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112270 48636
rect 119200 48384 119800 48496
rect 3042 48076 3052 48132
rect 3108 48076 3500 48132
rect 3556 48076 59276 48132
rect 59332 48076 59342 48132
rect 200 47796 800 47824
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 96626 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96910 47852
rect 200 47740 2044 47796
rect 2100 47740 2110 47796
rect 200 47712 800 47740
rect 119200 47124 119800 47152
rect 118066 47068 118076 47124
rect 118132 47068 119800 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 81266 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81550 47068
rect 111986 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112270 47068
rect 119200 47040 119800 47068
rect 200 46452 800 46480
rect 200 46396 1820 46452
rect 1876 46396 1886 46452
rect 200 46368 800 46396
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 96626 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96910 46284
rect 119200 45696 119800 45808
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 81266 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81550 45500
rect 111986 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112270 45500
rect 2146 45276 2156 45332
rect 2212 45276 4060 45332
rect 4116 45276 4126 45332
rect 200 45108 800 45136
rect 119200 45108 119800 45136
rect 200 45052 1932 45108
rect 1988 45052 2604 45108
rect 2660 45052 2670 45108
rect 118066 45052 118076 45108
rect 118132 45052 119800 45108
rect 200 45024 800 45052
rect 119200 45024 119800 45052
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 96626 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96910 44716
rect 200 44436 800 44464
rect 200 44380 1820 44436
rect 1876 44380 1886 44436
rect 200 44352 800 44380
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 81266 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81550 43932
rect 111986 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112270 43932
rect 119200 43764 119800 43792
rect 118066 43708 118076 43764
rect 118132 43708 119800 43764
rect 119200 43680 119800 43708
rect 200 43008 800 43120
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 96626 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96910 43148
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 81266 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81550 42364
rect 111986 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112270 42364
rect 119200 42336 119800 42448
rect 200 41748 800 41776
rect 200 41692 1820 41748
rect 1876 41692 1886 41748
rect 200 41664 800 41692
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 96626 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96910 41580
rect 119200 41076 119800 41104
rect 118066 41020 118076 41076
rect 118132 41020 119800 41076
rect 119200 40992 119800 41020
rect 2258 40908 2268 40964
rect 2324 40908 59388 40964
rect 59444 40908 59948 40964
rect 60004 40908 60014 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 81266 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81550 40796
rect 111986 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112270 40796
rect 200 40404 800 40432
rect 200 40348 1820 40404
rect 1876 40348 1886 40404
rect 200 40320 800 40348
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 96626 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96910 40012
rect 119200 39648 119800 39760
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 81266 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81550 39228
rect 111986 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112270 39228
rect 200 39060 800 39088
rect 200 39004 1820 39060
rect 1876 39004 1886 39060
rect 200 38976 800 39004
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 96626 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96910 38444
rect 119200 38388 119800 38416
rect 118066 38332 118076 38388
rect 118132 38332 119800 38388
rect 119200 38304 119800 38332
rect 200 37632 800 37744
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 81266 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81550 37660
rect 111986 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112270 37660
rect 119200 37632 119800 37744
rect 200 37044 800 37072
rect 200 36988 1820 37044
rect 1876 36988 1886 37044
rect 200 36960 800 36988
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 96626 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96910 36876
rect 119200 36372 119800 36400
rect 117730 36316 117740 36372
rect 117796 36316 119800 36372
rect 119200 36288 119800 36316
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 81266 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81550 36092
rect 111986 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112270 36092
rect 200 35700 800 35728
rect 200 35644 1820 35700
rect 1876 35644 1886 35700
rect 200 35616 800 35644
rect 60274 35532 60284 35588
rect 60340 35532 116284 35588
rect 116340 35532 116844 35588
rect 116900 35532 116910 35588
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 96626 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96910 35308
rect 119200 34944 119800 35056
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 81266 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81550 34524
rect 111986 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112270 34524
rect 200 34272 800 34384
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 96626 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96910 33740
rect 119200 33600 119800 33712
rect 200 33012 800 33040
rect 200 32956 1820 33012
rect 1876 32956 1886 33012
rect 200 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 81266 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81550 32956
rect 111986 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112270 32956
rect 119200 32256 119800 32368
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 96626 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96910 32172
rect 200 31584 800 31696
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 81266 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81550 31388
rect 111986 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112270 31388
rect 119200 30996 119800 31024
rect 118066 30940 118076 30996
rect 118132 30940 119800 30996
rect 119200 30912 119800 30940
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 96626 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96910 30604
rect 200 30240 800 30352
rect 119200 30240 119800 30352
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 81266 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81550 29820
rect 111986 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112270 29820
rect 200 29652 800 29680
rect 200 29596 1820 29652
rect 1876 29596 1886 29652
rect 200 29568 800 29596
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 96626 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96910 29036
rect 119200 28980 119800 29008
rect 118066 28924 118076 28980
rect 118132 28924 119800 28980
rect 119200 28896 119800 28924
rect 200 28224 800 28336
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 81266 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81550 28252
rect 111986 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112270 28252
rect 119200 27552 119800 27664
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 96626 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96910 27468
rect 200 26880 800 26992
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 81266 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81550 26684
rect 111986 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112270 26684
rect 119200 26292 119800 26320
rect 118066 26236 118076 26292
rect 118132 26236 119800 26292
rect 119200 26208 119800 26236
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 96626 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96910 25900
rect 200 25620 800 25648
rect 200 25564 1820 25620
rect 1876 25564 1886 25620
rect 200 25536 800 25564
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 81266 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81550 25116
rect 111986 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112270 25116
rect 119200 24948 119800 24976
rect 118066 24892 118076 24948
rect 118132 24892 119800 24948
rect 119200 24864 119800 24892
rect 200 24192 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 96626 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96910 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 81266 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81550 23548
rect 111986 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112270 23548
rect 119200 23520 119800 23632
rect 200 22932 800 22960
rect 119200 22932 119800 22960
rect 200 22876 1820 22932
rect 1876 22876 1886 22932
rect 118066 22876 118076 22932
rect 118132 22876 119800 22932
rect 200 22848 800 22876
rect 119200 22848 119800 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 96626 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96910 22764
rect 200 22176 800 22288
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 81266 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81550 21980
rect 111986 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112270 21980
rect 119200 21504 119800 21616
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 96626 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96910 21196
rect 200 20916 800 20944
rect 200 20860 1820 20916
rect 1876 20860 1886 20916
rect 200 20832 800 20860
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 81266 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81550 20412
rect 111986 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112270 20412
rect 119200 20244 119800 20272
rect 118066 20188 118076 20244
rect 118132 20188 119800 20244
rect 119200 20160 119800 20188
rect 200 19488 800 19600
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 96626 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96910 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 81266 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81550 18844
rect 111986 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112270 18844
rect 119200 18816 119800 18928
rect 200 18228 800 18256
rect 200 18172 1820 18228
rect 1876 18172 1886 18228
rect 200 18144 800 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 96626 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96910 18060
rect 119200 17556 119800 17584
rect 118066 17500 118076 17556
rect 118132 17500 119800 17556
rect 119200 17472 119800 17500
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 81266 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81550 17276
rect 111986 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112270 17276
rect 200 16884 800 16912
rect 200 16828 1820 16884
rect 1876 16828 1886 16884
rect 200 16800 800 16828
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 96626 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96910 16492
rect 119200 16212 119800 16240
rect 118066 16156 118076 16212
rect 118132 16156 119800 16212
rect 119200 16128 119800 16156
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 81266 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81550 15708
rect 111986 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112270 15708
rect 200 15456 800 15568
rect 119200 15456 119800 15568
rect 200 14784 800 14896
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 96626 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96910 14924
rect 119200 14196 119800 14224
rect 118066 14140 118076 14196
rect 118132 14140 119800 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 81266 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81550 14140
rect 111986 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112270 14140
rect 119200 14112 119800 14140
rect 200 13440 800 13552
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 96626 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96910 13356
rect 119200 12768 119800 12880
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 81266 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81550 12572
rect 111986 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112270 12572
rect 200 12096 800 12208
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 96626 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96910 11788
rect 119200 11508 119800 11536
rect 118066 11452 118076 11508
rect 118132 11452 119800 11508
rect 119200 11424 119800 11452
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 81266 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81550 11004
rect 111986 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112270 11004
rect 200 10836 800 10864
rect 200 10780 1820 10836
rect 1876 10780 1886 10836
rect 200 10752 800 10780
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 96626 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96910 10220
rect 119200 10164 119800 10192
rect 118066 10108 118076 10164
rect 118132 10108 119800 10164
rect 119200 10080 119800 10108
rect 200 9408 800 9520
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 81266 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81550 9436
rect 111986 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112270 9436
rect 119200 8736 119800 8848
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 96626 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96910 8652
rect 200 8064 800 8176
rect 119200 8064 119800 8176
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 81266 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81550 7868
rect 111986 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112270 7868
rect 200 7476 800 7504
rect 200 7420 1820 7476
rect 1876 7420 1886 7476
rect 200 7392 800 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 96626 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96910 7084
rect 119200 6720 119800 6832
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 81266 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81550 6300
rect 111986 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112270 6300
rect 200 6132 800 6160
rect 200 6076 1820 6132
rect 1876 6076 1886 6132
rect 200 6048 800 6076
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 96626 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96910 5516
rect 119200 5376 119800 5488
rect 200 4788 800 4816
rect 200 4732 1820 4788
rect 1876 4732 1886 4788
rect 200 4704 800 4732
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 81266 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81550 4732
rect 111986 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112270 4732
rect 20626 4172 20636 4228
rect 20692 4172 116508 4228
rect 116564 4172 116844 4228
rect 116900 4172 116910 4228
rect 119200 4116 119800 4144
rect 118066 4060 118076 4116
rect 118132 4060 119800 4116
rect 119200 4032 119800 4060
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 96626 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96910 3948
rect 200 3360 800 3472
rect 117730 3388 117740 3444
rect 117796 3388 119644 3444
rect 119700 3388 119710 3444
rect 68562 3276 68572 3332
rect 68628 3276 69132 3332
rect 69188 3276 69198 3332
rect 106866 3276 106876 3332
rect 106932 3276 107660 3332
rect 107716 3276 107726 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 81266 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81550 3164
rect 111986 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112270 3164
rect 119200 2688 119800 2800
rect 18 2268 28 2324
rect 84 2268 1820 2324
rect 1876 2268 1886 2324
rect 200 2016 800 2128
rect 119200 1344 119800 1456
rect 200 672 800 784
rect 119200 84 119800 112
rect 117954 28 117964 84
rect 118020 28 119800 84
rect 119200 0 119800 28
<< via3 >>
rect 4476 132468 4532 132524
rect 4580 132468 4636 132524
rect 4684 132468 4740 132524
rect 35196 132468 35252 132524
rect 35300 132468 35356 132524
rect 35404 132468 35460 132524
rect 65916 132468 65972 132524
rect 66020 132468 66076 132524
rect 66124 132468 66180 132524
rect 96636 132468 96692 132524
rect 96740 132468 96796 132524
rect 96844 132468 96900 132524
rect 19836 131684 19892 131740
rect 19940 131684 19996 131740
rect 20044 131684 20100 131740
rect 50556 131684 50612 131740
rect 50660 131684 50716 131740
rect 50764 131684 50820 131740
rect 81276 131684 81332 131740
rect 81380 131684 81436 131740
rect 81484 131684 81540 131740
rect 111996 131684 112052 131740
rect 112100 131684 112156 131740
rect 112204 131684 112260 131740
rect 4476 130900 4532 130956
rect 4580 130900 4636 130956
rect 4684 130900 4740 130956
rect 35196 130900 35252 130956
rect 35300 130900 35356 130956
rect 35404 130900 35460 130956
rect 65916 130900 65972 130956
rect 66020 130900 66076 130956
rect 66124 130900 66180 130956
rect 96636 130900 96692 130956
rect 96740 130900 96796 130956
rect 96844 130900 96900 130956
rect 19836 130116 19892 130172
rect 19940 130116 19996 130172
rect 20044 130116 20100 130172
rect 50556 130116 50612 130172
rect 50660 130116 50716 130172
rect 50764 130116 50820 130172
rect 81276 130116 81332 130172
rect 81380 130116 81436 130172
rect 81484 130116 81540 130172
rect 111996 130116 112052 130172
rect 112100 130116 112156 130172
rect 112204 130116 112260 130172
rect 4476 129332 4532 129388
rect 4580 129332 4636 129388
rect 4684 129332 4740 129388
rect 35196 129332 35252 129388
rect 35300 129332 35356 129388
rect 35404 129332 35460 129388
rect 65916 129332 65972 129388
rect 66020 129332 66076 129388
rect 66124 129332 66180 129388
rect 96636 129332 96692 129388
rect 96740 129332 96796 129388
rect 96844 129332 96900 129388
rect 19836 128548 19892 128604
rect 19940 128548 19996 128604
rect 20044 128548 20100 128604
rect 50556 128548 50612 128604
rect 50660 128548 50716 128604
rect 50764 128548 50820 128604
rect 81276 128548 81332 128604
rect 81380 128548 81436 128604
rect 81484 128548 81540 128604
rect 111996 128548 112052 128604
rect 112100 128548 112156 128604
rect 112204 128548 112260 128604
rect 4476 127764 4532 127820
rect 4580 127764 4636 127820
rect 4684 127764 4740 127820
rect 35196 127764 35252 127820
rect 35300 127764 35356 127820
rect 35404 127764 35460 127820
rect 65916 127764 65972 127820
rect 66020 127764 66076 127820
rect 66124 127764 66180 127820
rect 96636 127764 96692 127820
rect 96740 127764 96796 127820
rect 96844 127764 96900 127820
rect 19836 126980 19892 127036
rect 19940 126980 19996 127036
rect 20044 126980 20100 127036
rect 50556 126980 50612 127036
rect 50660 126980 50716 127036
rect 50764 126980 50820 127036
rect 81276 126980 81332 127036
rect 81380 126980 81436 127036
rect 81484 126980 81540 127036
rect 111996 126980 112052 127036
rect 112100 126980 112156 127036
rect 112204 126980 112260 127036
rect 4476 126196 4532 126252
rect 4580 126196 4636 126252
rect 4684 126196 4740 126252
rect 35196 126196 35252 126252
rect 35300 126196 35356 126252
rect 35404 126196 35460 126252
rect 65916 126196 65972 126252
rect 66020 126196 66076 126252
rect 66124 126196 66180 126252
rect 96636 126196 96692 126252
rect 96740 126196 96796 126252
rect 96844 126196 96900 126252
rect 19836 125412 19892 125468
rect 19940 125412 19996 125468
rect 20044 125412 20100 125468
rect 50556 125412 50612 125468
rect 50660 125412 50716 125468
rect 50764 125412 50820 125468
rect 81276 125412 81332 125468
rect 81380 125412 81436 125468
rect 81484 125412 81540 125468
rect 111996 125412 112052 125468
rect 112100 125412 112156 125468
rect 112204 125412 112260 125468
rect 4476 124628 4532 124684
rect 4580 124628 4636 124684
rect 4684 124628 4740 124684
rect 35196 124628 35252 124684
rect 35300 124628 35356 124684
rect 35404 124628 35460 124684
rect 65916 124628 65972 124684
rect 66020 124628 66076 124684
rect 66124 124628 66180 124684
rect 96636 124628 96692 124684
rect 96740 124628 96796 124684
rect 96844 124628 96900 124684
rect 19836 123844 19892 123900
rect 19940 123844 19996 123900
rect 20044 123844 20100 123900
rect 50556 123844 50612 123900
rect 50660 123844 50716 123900
rect 50764 123844 50820 123900
rect 81276 123844 81332 123900
rect 81380 123844 81436 123900
rect 81484 123844 81540 123900
rect 111996 123844 112052 123900
rect 112100 123844 112156 123900
rect 112204 123844 112260 123900
rect 4476 123060 4532 123116
rect 4580 123060 4636 123116
rect 4684 123060 4740 123116
rect 35196 123060 35252 123116
rect 35300 123060 35356 123116
rect 35404 123060 35460 123116
rect 65916 123060 65972 123116
rect 66020 123060 66076 123116
rect 66124 123060 66180 123116
rect 96636 123060 96692 123116
rect 96740 123060 96796 123116
rect 96844 123060 96900 123116
rect 19836 122276 19892 122332
rect 19940 122276 19996 122332
rect 20044 122276 20100 122332
rect 50556 122276 50612 122332
rect 50660 122276 50716 122332
rect 50764 122276 50820 122332
rect 81276 122276 81332 122332
rect 81380 122276 81436 122332
rect 81484 122276 81540 122332
rect 111996 122276 112052 122332
rect 112100 122276 112156 122332
rect 112204 122276 112260 122332
rect 4476 121492 4532 121548
rect 4580 121492 4636 121548
rect 4684 121492 4740 121548
rect 35196 121492 35252 121548
rect 35300 121492 35356 121548
rect 35404 121492 35460 121548
rect 65916 121492 65972 121548
rect 66020 121492 66076 121548
rect 66124 121492 66180 121548
rect 96636 121492 96692 121548
rect 96740 121492 96796 121548
rect 96844 121492 96900 121548
rect 19836 120708 19892 120764
rect 19940 120708 19996 120764
rect 20044 120708 20100 120764
rect 50556 120708 50612 120764
rect 50660 120708 50716 120764
rect 50764 120708 50820 120764
rect 81276 120708 81332 120764
rect 81380 120708 81436 120764
rect 81484 120708 81540 120764
rect 111996 120708 112052 120764
rect 112100 120708 112156 120764
rect 112204 120708 112260 120764
rect 4476 119924 4532 119980
rect 4580 119924 4636 119980
rect 4684 119924 4740 119980
rect 35196 119924 35252 119980
rect 35300 119924 35356 119980
rect 35404 119924 35460 119980
rect 65916 119924 65972 119980
rect 66020 119924 66076 119980
rect 66124 119924 66180 119980
rect 96636 119924 96692 119980
rect 96740 119924 96796 119980
rect 96844 119924 96900 119980
rect 19836 119140 19892 119196
rect 19940 119140 19996 119196
rect 20044 119140 20100 119196
rect 50556 119140 50612 119196
rect 50660 119140 50716 119196
rect 50764 119140 50820 119196
rect 81276 119140 81332 119196
rect 81380 119140 81436 119196
rect 81484 119140 81540 119196
rect 111996 119140 112052 119196
rect 112100 119140 112156 119196
rect 112204 119140 112260 119196
rect 4476 118356 4532 118412
rect 4580 118356 4636 118412
rect 4684 118356 4740 118412
rect 35196 118356 35252 118412
rect 35300 118356 35356 118412
rect 35404 118356 35460 118412
rect 65916 118356 65972 118412
rect 66020 118356 66076 118412
rect 66124 118356 66180 118412
rect 96636 118356 96692 118412
rect 96740 118356 96796 118412
rect 96844 118356 96900 118412
rect 19836 117572 19892 117628
rect 19940 117572 19996 117628
rect 20044 117572 20100 117628
rect 50556 117572 50612 117628
rect 50660 117572 50716 117628
rect 50764 117572 50820 117628
rect 81276 117572 81332 117628
rect 81380 117572 81436 117628
rect 81484 117572 81540 117628
rect 111996 117572 112052 117628
rect 112100 117572 112156 117628
rect 112204 117572 112260 117628
rect 4476 116788 4532 116844
rect 4580 116788 4636 116844
rect 4684 116788 4740 116844
rect 35196 116788 35252 116844
rect 35300 116788 35356 116844
rect 35404 116788 35460 116844
rect 65916 116788 65972 116844
rect 66020 116788 66076 116844
rect 66124 116788 66180 116844
rect 96636 116788 96692 116844
rect 96740 116788 96796 116844
rect 96844 116788 96900 116844
rect 19836 116004 19892 116060
rect 19940 116004 19996 116060
rect 20044 116004 20100 116060
rect 50556 116004 50612 116060
rect 50660 116004 50716 116060
rect 50764 116004 50820 116060
rect 81276 116004 81332 116060
rect 81380 116004 81436 116060
rect 81484 116004 81540 116060
rect 111996 116004 112052 116060
rect 112100 116004 112156 116060
rect 112204 116004 112260 116060
rect 4476 115220 4532 115276
rect 4580 115220 4636 115276
rect 4684 115220 4740 115276
rect 35196 115220 35252 115276
rect 35300 115220 35356 115276
rect 35404 115220 35460 115276
rect 65916 115220 65972 115276
rect 66020 115220 66076 115276
rect 66124 115220 66180 115276
rect 96636 115220 96692 115276
rect 96740 115220 96796 115276
rect 96844 115220 96900 115276
rect 19836 114436 19892 114492
rect 19940 114436 19996 114492
rect 20044 114436 20100 114492
rect 50556 114436 50612 114492
rect 50660 114436 50716 114492
rect 50764 114436 50820 114492
rect 81276 114436 81332 114492
rect 81380 114436 81436 114492
rect 81484 114436 81540 114492
rect 111996 114436 112052 114492
rect 112100 114436 112156 114492
rect 112204 114436 112260 114492
rect 4476 113652 4532 113708
rect 4580 113652 4636 113708
rect 4684 113652 4740 113708
rect 35196 113652 35252 113708
rect 35300 113652 35356 113708
rect 35404 113652 35460 113708
rect 65916 113652 65972 113708
rect 66020 113652 66076 113708
rect 66124 113652 66180 113708
rect 96636 113652 96692 113708
rect 96740 113652 96796 113708
rect 96844 113652 96900 113708
rect 19836 112868 19892 112924
rect 19940 112868 19996 112924
rect 20044 112868 20100 112924
rect 50556 112868 50612 112924
rect 50660 112868 50716 112924
rect 50764 112868 50820 112924
rect 81276 112868 81332 112924
rect 81380 112868 81436 112924
rect 81484 112868 81540 112924
rect 111996 112868 112052 112924
rect 112100 112868 112156 112924
rect 112204 112868 112260 112924
rect 4476 112084 4532 112140
rect 4580 112084 4636 112140
rect 4684 112084 4740 112140
rect 35196 112084 35252 112140
rect 35300 112084 35356 112140
rect 35404 112084 35460 112140
rect 65916 112084 65972 112140
rect 66020 112084 66076 112140
rect 66124 112084 66180 112140
rect 96636 112084 96692 112140
rect 96740 112084 96796 112140
rect 96844 112084 96900 112140
rect 19836 111300 19892 111356
rect 19940 111300 19996 111356
rect 20044 111300 20100 111356
rect 50556 111300 50612 111356
rect 50660 111300 50716 111356
rect 50764 111300 50820 111356
rect 81276 111300 81332 111356
rect 81380 111300 81436 111356
rect 81484 111300 81540 111356
rect 111996 111300 112052 111356
rect 112100 111300 112156 111356
rect 112204 111300 112260 111356
rect 4476 110516 4532 110572
rect 4580 110516 4636 110572
rect 4684 110516 4740 110572
rect 35196 110516 35252 110572
rect 35300 110516 35356 110572
rect 35404 110516 35460 110572
rect 65916 110516 65972 110572
rect 66020 110516 66076 110572
rect 66124 110516 66180 110572
rect 96636 110516 96692 110572
rect 96740 110516 96796 110572
rect 96844 110516 96900 110572
rect 19836 109732 19892 109788
rect 19940 109732 19996 109788
rect 20044 109732 20100 109788
rect 50556 109732 50612 109788
rect 50660 109732 50716 109788
rect 50764 109732 50820 109788
rect 81276 109732 81332 109788
rect 81380 109732 81436 109788
rect 81484 109732 81540 109788
rect 111996 109732 112052 109788
rect 112100 109732 112156 109788
rect 112204 109732 112260 109788
rect 4476 108948 4532 109004
rect 4580 108948 4636 109004
rect 4684 108948 4740 109004
rect 35196 108948 35252 109004
rect 35300 108948 35356 109004
rect 35404 108948 35460 109004
rect 65916 108948 65972 109004
rect 66020 108948 66076 109004
rect 66124 108948 66180 109004
rect 96636 108948 96692 109004
rect 96740 108948 96796 109004
rect 96844 108948 96900 109004
rect 19836 108164 19892 108220
rect 19940 108164 19996 108220
rect 20044 108164 20100 108220
rect 50556 108164 50612 108220
rect 50660 108164 50716 108220
rect 50764 108164 50820 108220
rect 81276 108164 81332 108220
rect 81380 108164 81436 108220
rect 81484 108164 81540 108220
rect 111996 108164 112052 108220
rect 112100 108164 112156 108220
rect 112204 108164 112260 108220
rect 4476 107380 4532 107436
rect 4580 107380 4636 107436
rect 4684 107380 4740 107436
rect 35196 107380 35252 107436
rect 35300 107380 35356 107436
rect 35404 107380 35460 107436
rect 65916 107380 65972 107436
rect 66020 107380 66076 107436
rect 66124 107380 66180 107436
rect 96636 107380 96692 107436
rect 96740 107380 96796 107436
rect 96844 107380 96900 107436
rect 19836 106596 19892 106652
rect 19940 106596 19996 106652
rect 20044 106596 20100 106652
rect 50556 106596 50612 106652
rect 50660 106596 50716 106652
rect 50764 106596 50820 106652
rect 81276 106596 81332 106652
rect 81380 106596 81436 106652
rect 81484 106596 81540 106652
rect 111996 106596 112052 106652
rect 112100 106596 112156 106652
rect 112204 106596 112260 106652
rect 4476 105812 4532 105868
rect 4580 105812 4636 105868
rect 4684 105812 4740 105868
rect 35196 105812 35252 105868
rect 35300 105812 35356 105868
rect 35404 105812 35460 105868
rect 65916 105812 65972 105868
rect 66020 105812 66076 105868
rect 66124 105812 66180 105868
rect 96636 105812 96692 105868
rect 96740 105812 96796 105868
rect 96844 105812 96900 105868
rect 19836 105028 19892 105084
rect 19940 105028 19996 105084
rect 20044 105028 20100 105084
rect 50556 105028 50612 105084
rect 50660 105028 50716 105084
rect 50764 105028 50820 105084
rect 81276 105028 81332 105084
rect 81380 105028 81436 105084
rect 81484 105028 81540 105084
rect 111996 105028 112052 105084
rect 112100 105028 112156 105084
rect 112204 105028 112260 105084
rect 4476 104244 4532 104300
rect 4580 104244 4636 104300
rect 4684 104244 4740 104300
rect 35196 104244 35252 104300
rect 35300 104244 35356 104300
rect 35404 104244 35460 104300
rect 65916 104244 65972 104300
rect 66020 104244 66076 104300
rect 66124 104244 66180 104300
rect 96636 104244 96692 104300
rect 96740 104244 96796 104300
rect 96844 104244 96900 104300
rect 19836 103460 19892 103516
rect 19940 103460 19996 103516
rect 20044 103460 20100 103516
rect 50556 103460 50612 103516
rect 50660 103460 50716 103516
rect 50764 103460 50820 103516
rect 81276 103460 81332 103516
rect 81380 103460 81436 103516
rect 81484 103460 81540 103516
rect 111996 103460 112052 103516
rect 112100 103460 112156 103516
rect 112204 103460 112260 103516
rect 4476 102676 4532 102732
rect 4580 102676 4636 102732
rect 4684 102676 4740 102732
rect 35196 102676 35252 102732
rect 35300 102676 35356 102732
rect 35404 102676 35460 102732
rect 65916 102676 65972 102732
rect 66020 102676 66076 102732
rect 66124 102676 66180 102732
rect 96636 102676 96692 102732
rect 96740 102676 96796 102732
rect 96844 102676 96900 102732
rect 19836 101892 19892 101948
rect 19940 101892 19996 101948
rect 20044 101892 20100 101948
rect 50556 101892 50612 101948
rect 50660 101892 50716 101948
rect 50764 101892 50820 101948
rect 81276 101892 81332 101948
rect 81380 101892 81436 101948
rect 81484 101892 81540 101948
rect 111996 101892 112052 101948
rect 112100 101892 112156 101948
rect 112204 101892 112260 101948
rect 4476 101108 4532 101164
rect 4580 101108 4636 101164
rect 4684 101108 4740 101164
rect 35196 101108 35252 101164
rect 35300 101108 35356 101164
rect 35404 101108 35460 101164
rect 65916 101108 65972 101164
rect 66020 101108 66076 101164
rect 66124 101108 66180 101164
rect 96636 101108 96692 101164
rect 96740 101108 96796 101164
rect 96844 101108 96900 101164
rect 19836 100324 19892 100380
rect 19940 100324 19996 100380
rect 20044 100324 20100 100380
rect 50556 100324 50612 100380
rect 50660 100324 50716 100380
rect 50764 100324 50820 100380
rect 81276 100324 81332 100380
rect 81380 100324 81436 100380
rect 81484 100324 81540 100380
rect 111996 100324 112052 100380
rect 112100 100324 112156 100380
rect 112204 100324 112260 100380
rect 4476 99540 4532 99596
rect 4580 99540 4636 99596
rect 4684 99540 4740 99596
rect 35196 99540 35252 99596
rect 35300 99540 35356 99596
rect 35404 99540 35460 99596
rect 65916 99540 65972 99596
rect 66020 99540 66076 99596
rect 66124 99540 66180 99596
rect 96636 99540 96692 99596
rect 96740 99540 96796 99596
rect 96844 99540 96900 99596
rect 19836 98756 19892 98812
rect 19940 98756 19996 98812
rect 20044 98756 20100 98812
rect 50556 98756 50612 98812
rect 50660 98756 50716 98812
rect 50764 98756 50820 98812
rect 81276 98756 81332 98812
rect 81380 98756 81436 98812
rect 81484 98756 81540 98812
rect 111996 98756 112052 98812
rect 112100 98756 112156 98812
rect 112204 98756 112260 98812
rect 4476 97972 4532 98028
rect 4580 97972 4636 98028
rect 4684 97972 4740 98028
rect 35196 97972 35252 98028
rect 35300 97972 35356 98028
rect 35404 97972 35460 98028
rect 65916 97972 65972 98028
rect 66020 97972 66076 98028
rect 66124 97972 66180 98028
rect 96636 97972 96692 98028
rect 96740 97972 96796 98028
rect 96844 97972 96900 98028
rect 19836 97188 19892 97244
rect 19940 97188 19996 97244
rect 20044 97188 20100 97244
rect 50556 97188 50612 97244
rect 50660 97188 50716 97244
rect 50764 97188 50820 97244
rect 81276 97188 81332 97244
rect 81380 97188 81436 97244
rect 81484 97188 81540 97244
rect 111996 97188 112052 97244
rect 112100 97188 112156 97244
rect 112204 97188 112260 97244
rect 4476 96404 4532 96460
rect 4580 96404 4636 96460
rect 4684 96404 4740 96460
rect 35196 96404 35252 96460
rect 35300 96404 35356 96460
rect 35404 96404 35460 96460
rect 65916 96404 65972 96460
rect 66020 96404 66076 96460
rect 66124 96404 66180 96460
rect 96636 96404 96692 96460
rect 96740 96404 96796 96460
rect 96844 96404 96900 96460
rect 19836 95620 19892 95676
rect 19940 95620 19996 95676
rect 20044 95620 20100 95676
rect 50556 95620 50612 95676
rect 50660 95620 50716 95676
rect 50764 95620 50820 95676
rect 81276 95620 81332 95676
rect 81380 95620 81436 95676
rect 81484 95620 81540 95676
rect 111996 95620 112052 95676
rect 112100 95620 112156 95676
rect 112204 95620 112260 95676
rect 4476 94836 4532 94892
rect 4580 94836 4636 94892
rect 4684 94836 4740 94892
rect 35196 94836 35252 94892
rect 35300 94836 35356 94892
rect 35404 94836 35460 94892
rect 65916 94836 65972 94892
rect 66020 94836 66076 94892
rect 66124 94836 66180 94892
rect 96636 94836 96692 94892
rect 96740 94836 96796 94892
rect 96844 94836 96900 94892
rect 19836 94052 19892 94108
rect 19940 94052 19996 94108
rect 20044 94052 20100 94108
rect 50556 94052 50612 94108
rect 50660 94052 50716 94108
rect 50764 94052 50820 94108
rect 81276 94052 81332 94108
rect 81380 94052 81436 94108
rect 81484 94052 81540 94108
rect 111996 94052 112052 94108
rect 112100 94052 112156 94108
rect 112204 94052 112260 94108
rect 4476 93268 4532 93324
rect 4580 93268 4636 93324
rect 4684 93268 4740 93324
rect 35196 93268 35252 93324
rect 35300 93268 35356 93324
rect 35404 93268 35460 93324
rect 65916 93268 65972 93324
rect 66020 93268 66076 93324
rect 66124 93268 66180 93324
rect 96636 93268 96692 93324
rect 96740 93268 96796 93324
rect 96844 93268 96900 93324
rect 19836 92484 19892 92540
rect 19940 92484 19996 92540
rect 20044 92484 20100 92540
rect 50556 92484 50612 92540
rect 50660 92484 50716 92540
rect 50764 92484 50820 92540
rect 81276 92484 81332 92540
rect 81380 92484 81436 92540
rect 81484 92484 81540 92540
rect 111996 92484 112052 92540
rect 112100 92484 112156 92540
rect 112204 92484 112260 92540
rect 4476 91700 4532 91756
rect 4580 91700 4636 91756
rect 4684 91700 4740 91756
rect 35196 91700 35252 91756
rect 35300 91700 35356 91756
rect 35404 91700 35460 91756
rect 65916 91700 65972 91756
rect 66020 91700 66076 91756
rect 66124 91700 66180 91756
rect 96636 91700 96692 91756
rect 96740 91700 96796 91756
rect 96844 91700 96900 91756
rect 19836 90916 19892 90972
rect 19940 90916 19996 90972
rect 20044 90916 20100 90972
rect 50556 90916 50612 90972
rect 50660 90916 50716 90972
rect 50764 90916 50820 90972
rect 81276 90916 81332 90972
rect 81380 90916 81436 90972
rect 81484 90916 81540 90972
rect 111996 90916 112052 90972
rect 112100 90916 112156 90972
rect 112204 90916 112260 90972
rect 4476 90132 4532 90188
rect 4580 90132 4636 90188
rect 4684 90132 4740 90188
rect 35196 90132 35252 90188
rect 35300 90132 35356 90188
rect 35404 90132 35460 90188
rect 65916 90132 65972 90188
rect 66020 90132 66076 90188
rect 66124 90132 66180 90188
rect 96636 90132 96692 90188
rect 96740 90132 96796 90188
rect 96844 90132 96900 90188
rect 19836 89348 19892 89404
rect 19940 89348 19996 89404
rect 20044 89348 20100 89404
rect 50556 89348 50612 89404
rect 50660 89348 50716 89404
rect 50764 89348 50820 89404
rect 81276 89348 81332 89404
rect 81380 89348 81436 89404
rect 81484 89348 81540 89404
rect 111996 89348 112052 89404
rect 112100 89348 112156 89404
rect 112204 89348 112260 89404
rect 4476 88564 4532 88620
rect 4580 88564 4636 88620
rect 4684 88564 4740 88620
rect 35196 88564 35252 88620
rect 35300 88564 35356 88620
rect 35404 88564 35460 88620
rect 65916 88564 65972 88620
rect 66020 88564 66076 88620
rect 66124 88564 66180 88620
rect 96636 88564 96692 88620
rect 96740 88564 96796 88620
rect 96844 88564 96900 88620
rect 19836 87780 19892 87836
rect 19940 87780 19996 87836
rect 20044 87780 20100 87836
rect 50556 87780 50612 87836
rect 50660 87780 50716 87836
rect 50764 87780 50820 87836
rect 81276 87780 81332 87836
rect 81380 87780 81436 87836
rect 81484 87780 81540 87836
rect 111996 87780 112052 87836
rect 112100 87780 112156 87836
rect 112204 87780 112260 87836
rect 4476 86996 4532 87052
rect 4580 86996 4636 87052
rect 4684 86996 4740 87052
rect 35196 86996 35252 87052
rect 35300 86996 35356 87052
rect 35404 86996 35460 87052
rect 65916 86996 65972 87052
rect 66020 86996 66076 87052
rect 66124 86996 66180 87052
rect 96636 86996 96692 87052
rect 96740 86996 96796 87052
rect 96844 86996 96900 87052
rect 19836 86212 19892 86268
rect 19940 86212 19996 86268
rect 20044 86212 20100 86268
rect 50556 86212 50612 86268
rect 50660 86212 50716 86268
rect 50764 86212 50820 86268
rect 81276 86212 81332 86268
rect 81380 86212 81436 86268
rect 81484 86212 81540 86268
rect 111996 86212 112052 86268
rect 112100 86212 112156 86268
rect 112204 86212 112260 86268
rect 4476 85428 4532 85484
rect 4580 85428 4636 85484
rect 4684 85428 4740 85484
rect 35196 85428 35252 85484
rect 35300 85428 35356 85484
rect 35404 85428 35460 85484
rect 65916 85428 65972 85484
rect 66020 85428 66076 85484
rect 66124 85428 66180 85484
rect 96636 85428 96692 85484
rect 96740 85428 96796 85484
rect 96844 85428 96900 85484
rect 19836 84644 19892 84700
rect 19940 84644 19996 84700
rect 20044 84644 20100 84700
rect 50556 84644 50612 84700
rect 50660 84644 50716 84700
rect 50764 84644 50820 84700
rect 81276 84644 81332 84700
rect 81380 84644 81436 84700
rect 81484 84644 81540 84700
rect 111996 84644 112052 84700
rect 112100 84644 112156 84700
rect 112204 84644 112260 84700
rect 4476 83860 4532 83916
rect 4580 83860 4636 83916
rect 4684 83860 4740 83916
rect 35196 83860 35252 83916
rect 35300 83860 35356 83916
rect 35404 83860 35460 83916
rect 65916 83860 65972 83916
rect 66020 83860 66076 83916
rect 66124 83860 66180 83916
rect 96636 83860 96692 83916
rect 96740 83860 96796 83916
rect 96844 83860 96900 83916
rect 19836 83076 19892 83132
rect 19940 83076 19996 83132
rect 20044 83076 20100 83132
rect 50556 83076 50612 83132
rect 50660 83076 50716 83132
rect 50764 83076 50820 83132
rect 81276 83076 81332 83132
rect 81380 83076 81436 83132
rect 81484 83076 81540 83132
rect 111996 83076 112052 83132
rect 112100 83076 112156 83132
rect 112204 83076 112260 83132
rect 4476 82292 4532 82348
rect 4580 82292 4636 82348
rect 4684 82292 4740 82348
rect 35196 82292 35252 82348
rect 35300 82292 35356 82348
rect 35404 82292 35460 82348
rect 65916 82292 65972 82348
rect 66020 82292 66076 82348
rect 66124 82292 66180 82348
rect 96636 82292 96692 82348
rect 96740 82292 96796 82348
rect 96844 82292 96900 82348
rect 19836 81508 19892 81564
rect 19940 81508 19996 81564
rect 20044 81508 20100 81564
rect 50556 81508 50612 81564
rect 50660 81508 50716 81564
rect 50764 81508 50820 81564
rect 81276 81508 81332 81564
rect 81380 81508 81436 81564
rect 81484 81508 81540 81564
rect 111996 81508 112052 81564
rect 112100 81508 112156 81564
rect 112204 81508 112260 81564
rect 4476 80724 4532 80780
rect 4580 80724 4636 80780
rect 4684 80724 4740 80780
rect 35196 80724 35252 80780
rect 35300 80724 35356 80780
rect 35404 80724 35460 80780
rect 65916 80724 65972 80780
rect 66020 80724 66076 80780
rect 66124 80724 66180 80780
rect 96636 80724 96692 80780
rect 96740 80724 96796 80780
rect 96844 80724 96900 80780
rect 19836 79940 19892 79996
rect 19940 79940 19996 79996
rect 20044 79940 20100 79996
rect 50556 79940 50612 79996
rect 50660 79940 50716 79996
rect 50764 79940 50820 79996
rect 81276 79940 81332 79996
rect 81380 79940 81436 79996
rect 81484 79940 81540 79996
rect 111996 79940 112052 79996
rect 112100 79940 112156 79996
rect 112204 79940 112260 79996
rect 4476 79156 4532 79212
rect 4580 79156 4636 79212
rect 4684 79156 4740 79212
rect 35196 79156 35252 79212
rect 35300 79156 35356 79212
rect 35404 79156 35460 79212
rect 65916 79156 65972 79212
rect 66020 79156 66076 79212
rect 66124 79156 66180 79212
rect 96636 79156 96692 79212
rect 96740 79156 96796 79212
rect 96844 79156 96900 79212
rect 19836 78372 19892 78428
rect 19940 78372 19996 78428
rect 20044 78372 20100 78428
rect 50556 78372 50612 78428
rect 50660 78372 50716 78428
rect 50764 78372 50820 78428
rect 81276 78372 81332 78428
rect 81380 78372 81436 78428
rect 81484 78372 81540 78428
rect 111996 78372 112052 78428
rect 112100 78372 112156 78428
rect 112204 78372 112260 78428
rect 4476 77588 4532 77644
rect 4580 77588 4636 77644
rect 4684 77588 4740 77644
rect 35196 77588 35252 77644
rect 35300 77588 35356 77644
rect 35404 77588 35460 77644
rect 65916 77588 65972 77644
rect 66020 77588 66076 77644
rect 66124 77588 66180 77644
rect 96636 77588 96692 77644
rect 96740 77588 96796 77644
rect 96844 77588 96900 77644
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 81276 76804 81332 76860
rect 81380 76804 81436 76860
rect 81484 76804 81540 76860
rect 111996 76804 112052 76860
rect 112100 76804 112156 76860
rect 112204 76804 112260 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 96636 76020 96692 76076
rect 96740 76020 96796 76076
rect 96844 76020 96900 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 81276 75236 81332 75292
rect 81380 75236 81436 75292
rect 81484 75236 81540 75292
rect 111996 75236 112052 75292
rect 112100 75236 112156 75292
rect 112204 75236 112260 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 96636 74452 96692 74508
rect 96740 74452 96796 74508
rect 96844 74452 96900 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 81276 73668 81332 73724
rect 81380 73668 81436 73724
rect 81484 73668 81540 73724
rect 111996 73668 112052 73724
rect 112100 73668 112156 73724
rect 112204 73668 112260 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 96636 72884 96692 72940
rect 96740 72884 96796 72940
rect 96844 72884 96900 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 81276 72100 81332 72156
rect 81380 72100 81436 72156
rect 81484 72100 81540 72156
rect 111996 72100 112052 72156
rect 112100 72100 112156 72156
rect 112204 72100 112260 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 96636 71316 96692 71372
rect 96740 71316 96796 71372
rect 96844 71316 96900 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 81276 70532 81332 70588
rect 81380 70532 81436 70588
rect 81484 70532 81540 70588
rect 111996 70532 112052 70588
rect 112100 70532 112156 70588
rect 112204 70532 112260 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 96636 69748 96692 69804
rect 96740 69748 96796 69804
rect 96844 69748 96900 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 81276 68964 81332 69020
rect 81380 68964 81436 69020
rect 81484 68964 81540 69020
rect 111996 68964 112052 69020
rect 112100 68964 112156 69020
rect 112204 68964 112260 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 96636 68180 96692 68236
rect 96740 68180 96796 68236
rect 96844 68180 96900 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 81276 67396 81332 67452
rect 81380 67396 81436 67452
rect 81484 67396 81540 67452
rect 111996 67396 112052 67452
rect 112100 67396 112156 67452
rect 112204 67396 112260 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 96636 66612 96692 66668
rect 96740 66612 96796 66668
rect 96844 66612 96900 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 81276 65828 81332 65884
rect 81380 65828 81436 65884
rect 81484 65828 81540 65884
rect 111996 65828 112052 65884
rect 112100 65828 112156 65884
rect 112204 65828 112260 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 96636 65044 96692 65100
rect 96740 65044 96796 65100
rect 96844 65044 96900 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 81276 64260 81332 64316
rect 81380 64260 81436 64316
rect 81484 64260 81540 64316
rect 111996 64260 112052 64316
rect 112100 64260 112156 64316
rect 112204 64260 112260 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 96636 63476 96692 63532
rect 96740 63476 96796 63532
rect 96844 63476 96900 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 81276 62692 81332 62748
rect 81380 62692 81436 62748
rect 81484 62692 81540 62748
rect 111996 62692 112052 62748
rect 112100 62692 112156 62748
rect 112204 62692 112260 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 96636 61908 96692 61964
rect 96740 61908 96796 61964
rect 96844 61908 96900 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 81276 61124 81332 61180
rect 81380 61124 81436 61180
rect 81484 61124 81540 61180
rect 111996 61124 112052 61180
rect 112100 61124 112156 61180
rect 112204 61124 112260 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 96636 60340 96692 60396
rect 96740 60340 96796 60396
rect 96844 60340 96900 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 81276 59556 81332 59612
rect 81380 59556 81436 59612
rect 81484 59556 81540 59612
rect 111996 59556 112052 59612
rect 112100 59556 112156 59612
rect 112204 59556 112260 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 96636 58772 96692 58828
rect 96740 58772 96796 58828
rect 96844 58772 96900 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 81276 57988 81332 58044
rect 81380 57988 81436 58044
rect 81484 57988 81540 58044
rect 111996 57988 112052 58044
rect 112100 57988 112156 58044
rect 112204 57988 112260 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 96636 57204 96692 57260
rect 96740 57204 96796 57260
rect 96844 57204 96900 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 81276 56420 81332 56476
rect 81380 56420 81436 56476
rect 81484 56420 81540 56476
rect 111996 56420 112052 56476
rect 112100 56420 112156 56476
rect 112204 56420 112260 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 96636 55636 96692 55692
rect 96740 55636 96796 55692
rect 96844 55636 96900 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 81276 54852 81332 54908
rect 81380 54852 81436 54908
rect 81484 54852 81540 54908
rect 111996 54852 112052 54908
rect 112100 54852 112156 54908
rect 112204 54852 112260 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 96636 54068 96692 54124
rect 96740 54068 96796 54124
rect 96844 54068 96900 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 81276 53284 81332 53340
rect 81380 53284 81436 53340
rect 81484 53284 81540 53340
rect 111996 53284 112052 53340
rect 112100 53284 112156 53340
rect 112204 53284 112260 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 96636 52500 96692 52556
rect 96740 52500 96796 52556
rect 96844 52500 96900 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 81276 51716 81332 51772
rect 81380 51716 81436 51772
rect 81484 51716 81540 51772
rect 111996 51716 112052 51772
rect 112100 51716 112156 51772
rect 112204 51716 112260 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 96636 50932 96692 50988
rect 96740 50932 96796 50988
rect 96844 50932 96900 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 81276 50148 81332 50204
rect 81380 50148 81436 50204
rect 81484 50148 81540 50204
rect 111996 50148 112052 50204
rect 112100 50148 112156 50204
rect 112204 50148 112260 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 96636 49364 96692 49420
rect 96740 49364 96796 49420
rect 96844 49364 96900 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 81276 48580 81332 48636
rect 81380 48580 81436 48636
rect 81484 48580 81540 48636
rect 111996 48580 112052 48636
rect 112100 48580 112156 48636
rect 112204 48580 112260 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 96636 47796 96692 47852
rect 96740 47796 96796 47852
rect 96844 47796 96900 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 81276 47012 81332 47068
rect 81380 47012 81436 47068
rect 81484 47012 81540 47068
rect 111996 47012 112052 47068
rect 112100 47012 112156 47068
rect 112204 47012 112260 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 96636 46228 96692 46284
rect 96740 46228 96796 46284
rect 96844 46228 96900 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 81276 45444 81332 45500
rect 81380 45444 81436 45500
rect 81484 45444 81540 45500
rect 111996 45444 112052 45500
rect 112100 45444 112156 45500
rect 112204 45444 112260 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 96636 44660 96692 44716
rect 96740 44660 96796 44716
rect 96844 44660 96900 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 81276 43876 81332 43932
rect 81380 43876 81436 43932
rect 81484 43876 81540 43932
rect 111996 43876 112052 43932
rect 112100 43876 112156 43932
rect 112204 43876 112260 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 96636 43092 96692 43148
rect 96740 43092 96796 43148
rect 96844 43092 96900 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 81276 42308 81332 42364
rect 81380 42308 81436 42364
rect 81484 42308 81540 42364
rect 111996 42308 112052 42364
rect 112100 42308 112156 42364
rect 112204 42308 112260 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 96636 41524 96692 41580
rect 96740 41524 96796 41580
rect 96844 41524 96900 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 81276 40740 81332 40796
rect 81380 40740 81436 40796
rect 81484 40740 81540 40796
rect 111996 40740 112052 40796
rect 112100 40740 112156 40796
rect 112204 40740 112260 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 96636 39956 96692 40012
rect 96740 39956 96796 40012
rect 96844 39956 96900 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 81276 39172 81332 39228
rect 81380 39172 81436 39228
rect 81484 39172 81540 39228
rect 111996 39172 112052 39228
rect 112100 39172 112156 39228
rect 112204 39172 112260 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 96636 38388 96692 38444
rect 96740 38388 96796 38444
rect 96844 38388 96900 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 81276 37604 81332 37660
rect 81380 37604 81436 37660
rect 81484 37604 81540 37660
rect 111996 37604 112052 37660
rect 112100 37604 112156 37660
rect 112204 37604 112260 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 96636 36820 96692 36876
rect 96740 36820 96796 36876
rect 96844 36820 96900 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 81276 36036 81332 36092
rect 81380 36036 81436 36092
rect 81484 36036 81540 36092
rect 111996 36036 112052 36092
rect 112100 36036 112156 36092
rect 112204 36036 112260 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 96636 35252 96692 35308
rect 96740 35252 96796 35308
rect 96844 35252 96900 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 81276 34468 81332 34524
rect 81380 34468 81436 34524
rect 81484 34468 81540 34524
rect 111996 34468 112052 34524
rect 112100 34468 112156 34524
rect 112204 34468 112260 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 96636 33684 96692 33740
rect 96740 33684 96796 33740
rect 96844 33684 96900 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 81276 32900 81332 32956
rect 81380 32900 81436 32956
rect 81484 32900 81540 32956
rect 111996 32900 112052 32956
rect 112100 32900 112156 32956
rect 112204 32900 112260 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 96636 32116 96692 32172
rect 96740 32116 96796 32172
rect 96844 32116 96900 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 81276 31332 81332 31388
rect 81380 31332 81436 31388
rect 81484 31332 81540 31388
rect 111996 31332 112052 31388
rect 112100 31332 112156 31388
rect 112204 31332 112260 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 96636 30548 96692 30604
rect 96740 30548 96796 30604
rect 96844 30548 96900 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 81276 29764 81332 29820
rect 81380 29764 81436 29820
rect 81484 29764 81540 29820
rect 111996 29764 112052 29820
rect 112100 29764 112156 29820
rect 112204 29764 112260 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 96636 28980 96692 29036
rect 96740 28980 96796 29036
rect 96844 28980 96900 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 81276 28196 81332 28252
rect 81380 28196 81436 28252
rect 81484 28196 81540 28252
rect 111996 28196 112052 28252
rect 112100 28196 112156 28252
rect 112204 28196 112260 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 96636 27412 96692 27468
rect 96740 27412 96796 27468
rect 96844 27412 96900 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 81276 26628 81332 26684
rect 81380 26628 81436 26684
rect 81484 26628 81540 26684
rect 111996 26628 112052 26684
rect 112100 26628 112156 26684
rect 112204 26628 112260 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 96636 25844 96692 25900
rect 96740 25844 96796 25900
rect 96844 25844 96900 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 81276 25060 81332 25116
rect 81380 25060 81436 25116
rect 81484 25060 81540 25116
rect 111996 25060 112052 25116
rect 112100 25060 112156 25116
rect 112204 25060 112260 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 96636 24276 96692 24332
rect 96740 24276 96796 24332
rect 96844 24276 96900 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 81276 23492 81332 23548
rect 81380 23492 81436 23548
rect 81484 23492 81540 23548
rect 111996 23492 112052 23548
rect 112100 23492 112156 23548
rect 112204 23492 112260 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 96636 22708 96692 22764
rect 96740 22708 96796 22764
rect 96844 22708 96900 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 81276 21924 81332 21980
rect 81380 21924 81436 21980
rect 81484 21924 81540 21980
rect 111996 21924 112052 21980
rect 112100 21924 112156 21980
rect 112204 21924 112260 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 96636 21140 96692 21196
rect 96740 21140 96796 21196
rect 96844 21140 96900 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 81276 20356 81332 20412
rect 81380 20356 81436 20412
rect 81484 20356 81540 20412
rect 111996 20356 112052 20412
rect 112100 20356 112156 20412
rect 112204 20356 112260 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 96636 19572 96692 19628
rect 96740 19572 96796 19628
rect 96844 19572 96900 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 81276 18788 81332 18844
rect 81380 18788 81436 18844
rect 81484 18788 81540 18844
rect 111996 18788 112052 18844
rect 112100 18788 112156 18844
rect 112204 18788 112260 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 96636 18004 96692 18060
rect 96740 18004 96796 18060
rect 96844 18004 96900 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 81276 17220 81332 17276
rect 81380 17220 81436 17276
rect 81484 17220 81540 17276
rect 111996 17220 112052 17276
rect 112100 17220 112156 17276
rect 112204 17220 112260 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 96636 16436 96692 16492
rect 96740 16436 96796 16492
rect 96844 16436 96900 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 81276 15652 81332 15708
rect 81380 15652 81436 15708
rect 81484 15652 81540 15708
rect 111996 15652 112052 15708
rect 112100 15652 112156 15708
rect 112204 15652 112260 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 96636 14868 96692 14924
rect 96740 14868 96796 14924
rect 96844 14868 96900 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 81276 14084 81332 14140
rect 81380 14084 81436 14140
rect 81484 14084 81540 14140
rect 111996 14084 112052 14140
rect 112100 14084 112156 14140
rect 112204 14084 112260 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 96636 13300 96692 13356
rect 96740 13300 96796 13356
rect 96844 13300 96900 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 81276 12516 81332 12572
rect 81380 12516 81436 12572
rect 81484 12516 81540 12572
rect 111996 12516 112052 12572
rect 112100 12516 112156 12572
rect 112204 12516 112260 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 96636 11732 96692 11788
rect 96740 11732 96796 11788
rect 96844 11732 96900 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 81276 10948 81332 11004
rect 81380 10948 81436 11004
rect 81484 10948 81540 11004
rect 111996 10948 112052 11004
rect 112100 10948 112156 11004
rect 112204 10948 112260 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 96636 10164 96692 10220
rect 96740 10164 96796 10220
rect 96844 10164 96900 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 81276 9380 81332 9436
rect 81380 9380 81436 9436
rect 81484 9380 81540 9436
rect 111996 9380 112052 9436
rect 112100 9380 112156 9436
rect 112204 9380 112260 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 96636 8596 96692 8652
rect 96740 8596 96796 8652
rect 96844 8596 96900 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 81276 7812 81332 7868
rect 81380 7812 81436 7868
rect 81484 7812 81540 7868
rect 111996 7812 112052 7868
rect 112100 7812 112156 7868
rect 112204 7812 112260 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 96636 7028 96692 7084
rect 96740 7028 96796 7084
rect 96844 7028 96900 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 81276 6244 81332 6300
rect 81380 6244 81436 6300
rect 81484 6244 81540 6300
rect 111996 6244 112052 6300
rect 112100 6244 112156 6300
rect 112204 6244 112260 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 96636 5460 96692 5516
rect 96740 5460 96796 5516
rect 96844 5460 96900 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 81276 4676 81332 4732
rect 81380 4676 81436 4732
rect 81484 4676 81540 4732
rect 111996 4676 112052 4732
rect 112100 4676 112156 4732
rect 112204 4676 112260 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 96636 3892 96692 3948
rect 96740 3892 96796 3948
rect 96844 3892 96900 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 81276 3108 81332 3164
rect 81380 3108 81436 3164
rect 81484 3108 81540 3164
rect 111996 3108 112052 3164
rect 112100 3108 112156 3164
rect 112204 3108 112260 3164
<< metal4 >>
rect 4448 132524 4768 132556
rect 4448 132468 4476 132524
rect 4532 132468 4580 132524
rect 4636 132468 4684 132524
rect 4740 132468 4768 132524
rect 4448 130956 4768 132468
rect 4448 130900 4476 130956
rect 4532 130900 4580 130956
rect 4636 130900 4684 130956
rect 4740 130900 4768 130956
rect 4448 129388 4768 130900
rect 4448 129332 4476 129388
rect 4532 129332 4580 129388
rect 4636 129332 4684 129388
rect 4740 129332 4768 129388
rect 4448 127820 4768 129332
rect 4448 127764 4476 127820
rect 4532 127764 4580 127820
rect 4636 127764 4684 127820
rect 4740 127764 4768 127820
rect 4448 126252 4768 127764
rect 4448 126196 4476 126252
rect 4532 126196 4580 126252
rect 4636 126196 4684 126252
rect 4740 126196 4768 126252
rect 4448 124684 4768 126196
rect 4448 124628 4476 124684
rect 4532 124628 4580 124684
rect 4636 124628 4684 124684
rect 4740 124628 4768 124684
rect 4448 123116 4768 124628
rect 4448 123060 4476 123116
rect 4532 123060 4580 123116
rect 4636 123060 4684 123116
rect 4740 123060 4768 123116
rect 4448 121548 4768 123060
rect 4448 121492 4476 121548
rect 4532 121492 4580 121548
rect 4636 121492 4684 121548
rect 4740 121492 4768 121548
rect 4448 119980 4768 121492
rect 4448 119924 4476 119980
rect 4532 119924 4580 119980
rect 4636 119924 4684 119980
rect 4740 119924 4768 119980
rect 4448 118412 4768 119924
rect 4448 118356 4476 118412
rect 4532 118356 4580 118412
rect 4636 118356 4684 118412
rect 4740 118356 4768 118412
rect 4448 116844 4768 118356
rect 4448 116788 4476 116844
rect 4532 116788 4580 116844
rect 4636 116788 4684 116844
rect 4740 116788 4768 116844
rect 4448 115276 4768 116788
rect 4448 115220 4476 115276
rect 4532 115220 4580 115276
rect 4636 115220 4684 115276
rect 4740 115220 4768 115276
rect 4448 113708 4768 115220
rect 4448 113652 4476 113708
rect 4532 113652 4580 113708
rect 4636 113652 4684 113708
rect 4740 113652 4768 113708
rect 4448 112140 4768 113652
rect 4448 112084 4476 112140
rect 4532 112084 4580 112140
rect 4636 112084 4684 112140
rect 4740 112084 4768 112140
rect 4448 110572 4768 112084
rect 4448 110516 4476 110572
rect 4532 110516 4580 110572
rect 4636 110516 4684 110572
rect 4740 110516 4768 110572
rect 4448 109004 4768 110516
rect 4448 108948 4476 109004
rect 4532 108948 4580 109004
rect 4636 108948 4684 109004
rect 4740 108948 4768 109004
rect 4448 107436 4768 108948
rect 4448 107380 4476 107436
rect 4532 107380 4580 107436
rect 4636 107380 4684 107436
rect 4740 107380 4768 107436
rect 4448 105868 4768 107380
rect 4448 105812 4476 105868
rect 4532 105812 4580 105868
rect 4636 105812 4684 105868
rect 4740 105812 4768 105868
rect 4448 104300 4768 105812
rect 4448 104244 4476 104300
rect 4532 104244 4580 104300
rect 4636 104244 4684 104300
rect 4740 104244 4768 104300
rect 4448 102732 4768 104244
rect 4448 102676 4476 102732
rect 4532 102676 4580 102732
rect 4636 102676 4684 102732
rect 4740 102676 4768 102732
rect 4448 101164 4768 102676
rect 4448 101108 4476 101164
rect 4532 101108 4580 101164
rect 4636 101108 4684 101164
rect 4740 101108 4768 101164
rect 4448 99596 4768 101108
rect 4448 99540 4476 99596
rect 4532 99540 4580 99596
rect 4636 99540 4684 99596
rect 4740 99540 4768 99596
rect 4448 98028 4768 99540
rect 4448 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4768 98028
rect 4448 96460 4768 97972
rect 4448 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4768 96460
rect 4448 94892 4768 96404
rect 4448 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4768 94892
rect 4448 93324 4768 94836
rect 4448 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4768 93324
rect 4448 91756 4768 93268
rect 4448 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4768 91756
rect 4448 90188 4768 91700
rect 4448 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4768 90188
rect 4448 88620 4768 90132
rect 4448 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4768 88620
rect 4448 87052 4768 88564
rect 4448 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4768 87052
rect 4448 85484 4768 86996
rect 4448 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4768 85484
rect 4448 83916 4768 85428
rect 4448 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4768 83916
rect 4448 82348 4768 83860
rect 4448 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4768 82348
rect 4448 80780 4768 82292
rect 4448 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4768 80780
rect 4448 79212 4768 80724
rect 4448 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4768 79212
rect 4448 77644 4768 79156
rect 4448 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4768 77644
rect 4448 76076 4768 77588
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 131740 20128 132556
rect 19808 131684 19836 131740
rect 19892 131684 19940 131740
rect 19996 131684 20044 131740
rect 20100 131684 20128 131740
rect 19808 130172 20128 131684
rect 19808 130116 19836 130172
rect 19892 130116 19940 130172
rect 19996 130116 20044 130172
rect 20100 130116 20128 130172
rect 19808 128604 20128 130116
rect 19808 128548 19836 128604
rect 19892 128548 19940 128604
rect 19996 128548 20044 128604
rect 20100 128548 20128 128604
rect 19808 127036 20128 128548
rect 19808 126980 19836 127036
rect 19892 126980 19940 127036
rect 19996 126980 20044 127036
rect 20100 126980 20128 127036
rect 19808 125468 20128 126980
rect 19808 125412 19836 125468
rect 19892 125412 19940 125468
rect 19996 125412 20044 125468
rect 20100 125412 20128 125468
rect 19808 123900 20128 125412
rect 19808 123844 19836 123900
rect 19892 123844 19940 123900
rect 19996 123844 20044 123900
rect 20100 123844 20128 123900
rect 19808 122332 20128 123844
rect 19808 122276 19836 122332
rect 19892 122276 19940 122332
rect 19996 122276 20044 122332
rect 20100 122276 20128 122332
rect 19808 120764 20128 122276
rect 19808 120708 19836 120764
rect 19892 120708 19940 120764
rect 19996 120708 20044 120764
rect 20100 120708 20128 120764
rect 19808 119196 20128 120708
rect 19808 119140 19836 119196
rect 19892 119140 19940 119196
rect 19996 119140 20044 119196
rect 20100 119140 20128 119196
rect 19808 117628 20128 119140
rect 19808 117572 19836 117628
rect 19892 117572 19940 117628
rect 19996 117572 20044 117628
rect 20100 117572 20128 117628
rect 19808 116060 20128 117572
rect 19808 116004 19836 116060
rect 19892 116004 19940 116060
rect 19996 116004 20044 116060
rect 20100 116004 20128 116060
rect 19808 114492 20128 116004
rect 19808 114436 19836 114492
rect 19892 114436 19940 114492
rect 19996 114436 20044 114492
rect 20100 114436 20128 114492
rect 19808 112924 20128 114436
rect 19808 112868 19836 112924
rect 19892 112868 19940 112924
rect 19996 112868 20044 112924
rect 20100 112868 20128 112924
rect 19808 111356 20128 112868
rect 19808 111300 19836 111356
rect 19892 111300 19940 111356
rect 19996 111300 20044 111356
rect 20100 111300 20128 111356
rect 19808 109788 20128 111300
rect 19808 109732 19836 109788
rect 19892 109732 19940 109788
rect 19996 109732 20044 109788
rect 20100 109732 20128 109788
rect 19808 108220 20128 109732
rect 19808 108164 19836 108220
rect 19892 108164 19940 108220
rect 19996 108164 20044 108220
rect 20100 108164 20128 108220
rect 19808 106652 20128 108164
rect 19808 106596 19836 106652
rect 19892 106596 19940 106652
rect 19996 106596 20044 106652
rect 20100 106596 20128 106652
rect 19808 105084 20128 106596
rect 19808 105028 19836 105084
rect 19892 105028 19940 105084
rect 19996 105028 20044 105084
rect 20100 105028 20128 105084
rect 19808 103516 20128 105028
rect 19808 103460 19836 103516
rect 19892 103460 19940 103516
rect 19996 103460 20044 103516
rect 20100 103460 20128 103516
rect 19808 101948 20128 103460
rect 19808 101892 19836 101948
rect 19892 101892 19940 101948
rect 19996 101892 20044 101948
rect 20100 101892 20128 101948
rect 19808 100380 20128 101892
rect 19808 100324 19836 100380
rect 19892 100324 19940 100380
rect 19996 100324 20044 100380
rect 20100 100324 20128 100380
rect 19808 98812 20128 100324
rect 19808 98756 19836 98812
rect 19892 98756 19940 98812
rect 19996 98756 20044 98812
rect 20100 98756 20128 98812
rect 19808 97244 20128 98756
rect 19808 97188 19836 97244
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 20100 97188 20128 97244
rect 19808 95676 20128 97188
rect 19808 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20128 95676
rect 19808 94108 20128 95620
rect 19808 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20128 94108
rect 19808 92540 20128 94052
rect 19808 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20128 92540
rect 19808 90972 20128 92484
rect 19808 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20128 90972
rect 19808 89404 20128 90916
rect 19808 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20128 89404
rect 19808 87836 20128 89348
rect 19808 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20128 87836
rect 19808 86268 20128 87780
rect 19808 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20128 86268
rect 19808 84700 20128 86212
rect 19808 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20128 84700
rect 19808 83132 20128 84644
rect 19808 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20128 83132
rect 19808 81564 20128 83076
rect 19808 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20128 81564
rect 19808 79996 20128 81508
rect 19808 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20128 79996
rect 19808 78428 20128 79940
rect 19808 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20128 78428
rect 19808 76860 20128 78372
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 132524 35488 132556
rect 35168 132468 35196 132524
rect 35252 132468 35300 132524
rect 35356 132468 35404 132524
rect 35460 132468 35488 132524
rect 35168 130956 35488 132468
rect 35168 130900 35196 130956
rect 35252 130900 35300 130956
rect 35356 130900 35404 130956
rect 35460 130900 35488 130956
rect 35168 129388 35488 130900
rect 35168 129332 35196 129388
rect 35252 129332 35300 129388
rect 35356 129332 35404 129388
rect 35460 129332 35488 129388
rect 35168 127820 35488 129332
rect 35168 127764 35196 127820
rect 35252 127764 35300 127820
rect 35356 127764 35404 127820
rect 35460 127764 35488 127820
rect 35168 126252 35488 127764
rect 35168 126196 35196 126252
rect 35252 126196 35300 126252
rect 35356 126196 35404 126252
rect 35460 126196 35488 126252
rect 35168 124684 35488 126196
rect 35168 124628 35196 124684
rect 35252 124628 35300 124684
rect 35356 124628 35404 124684
rect 35460 124628 35488 124684
rect 35168 123116 35488 124628
rect 35168 123060 35196 123116
rect 35252 123060 35300 123116
rect 35356 123060 35404 123116
rect 35460 123060 35488 123116
rect 35168 121548 35488 123060
rect 35168 121492 35196 121548
rect 35252 121492 35300 121548
rect 35356 121492 35404 121548
rect 35460 121492 35488 121548
rect 35168 119980 35488 121492
rect 35168 119924 35196 119980
rect 35252 119924 35300 119980
rect 35356 119924 35404 119980
rect 35460 119924 35488 119980
rect 35168 118412 35488 119924
rect 35168 118356 35196 118412
rect 35252 118356 35300 118412
rect 35356 118356 35404 118412
rect 35460 118356 35488 118412
rect 35168 116844 35488 118356
rect 35168 116788 35196 116844
rect 35252 116788 35300 116844
rect 35356 116788 35404 116844
rect 35460 116788 35488 116844
rect 35168 115276 35488 116788
rect 35168 115220 35196 115276
rect 35252 115220 35300 115276
rect 35356 115220 35404 115276
rect 35460 115220 35488 115276
rect 35168 113708 35488 115220
rect 35168 113652 35196 113708
rect 35252 113652 35300 113708
rect 35356 113652 35404 113708
rect 35460 113652 35488 113708
rect 35168 112140 35488 113652
rect 35168 112084 35196 112140
rect 35252 112084 35300 112140
rect 35356 112084 35404 112140
rect 35460 112084 35488 112140
rect 35168 110572 35488 112084
rect 35168 110516 35196 110572
rect 35252 110516 35300 110572
rect 35356 110516 35404 110572
rect 35460 110516 35488 110572
rect 35168 109004 35488 110516
rect 35168 108948 35196 109004
rect 35252 108948 35300 109004
rect 35356 108948 35404 109004
rect 35460 108948 35488 109004
rect 35168 107436 35488 108948
rect 35168 107380 35196 107436
rect 35252 107380 35300 107436
rect 35356 107380 35404 107436
rect 35460 107380 35488 107436
rect 35168 105868 35488 107380
rect 35168 105812 35196 105868
rect 35252 105812 35300 105868
rect 35356 105812 35404 105868
rect 35460 105812 35488 105868
rect 35168 104300 35488 105812
rect 35168 104244 35196 104300
rect 35252 104244 35300 104300
rect 35356 104244 35404 104300
rect 35460 104244 35488 104300
rect 35168 102732 35488 104244
rect 35168 102676 35196 102732
rect 35252 102676 35300 102732
rect 35356 102676 35404 102732
rect 35460 102676 35488 102732
rect 35168 101164 35488 102676
rect 35168 101108 35196 101164
rect 35252 101108 35300 101164
rect 35356 101108 35404 101164
rect 35460 101108 35488 101164
rect 35168 99596 35488 101108
rect 35168 99540 35196 99596
rect 35252 99540 35300 99596
rect 35356 99540 35404 99596
rect 35460 99540 35488 99596
rect 35168 98028 35488 99540
rect 35168 97972 35196 98028
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35460 97972 35488 98028
rect 35168 96460 35488 97972
rect 35168 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35488 96460
rect 35168 94892 35488 96404
rect 35168 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35488 94892
rect 35168 93324 35488 94836
rect 35168 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35488 93324
rect 35168 91756 35488 93268
rect 35168 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35488 91756
rect 35168 90188 35488 91700
rect 35168 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35488 90188
rect 35168 88620 35488 90132
rect 35168 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35488 88620
rect 35168 87052 35488 88564
rect 35168 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35488 87052
rect 35168 85484 35488 86996
rect 35168 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35488 85484
rect 35168 83916 35488 85428
rect 35168 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35488 83916
rect 35168 82348 35488 83860
rect 35168 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35488 82348
rect 35168 80780 35488 82292
rect 35168 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35488 80780
rect 35168 79212 35488 80724
rect 35168 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35488 79212
rect 35168 77644 35488 79156
rect 35168 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35488 77644
rect 35168 76076 35488 77588
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 131740 50848 132556
rect 50528 131684 50556 131740
rect 50612 131684 50660 131740
rect 50716 131684 50764 131740
rect 50820 131684 50848 131740
rect 50528 130172 50848 131684
rect 50528 130116 50556 130172
rect 50612 130116 50660 130172
rect 50716 130116 50764 130172
rect 50820 130116 50848 130172
rect 50528 128604 50848 130116
rect 50528 128548 50556 128604
rect 50612 128548 50660 128604
rect 50716 128548 50764 128604
rect 50820 128548 50848 128604
rect 50528 127036 50848 128548
rect 50528 126980 50556 127036
rect 50612 126980 50660 127036
rect 50716 126980 50764 127036
rect 50820 126980 50848 127036
rect 50528 125468 50848 126980
rect 50528 125412 50556 125468
rect 50612 125412 50660 125468
rect 50716 125412 50764 125468
rect 50820 125412 50848 125468
rect 50528 123900 50848 125412
rect 50528 123844 50556 123900
rect 50612 123844 50660 123900
rect 50716 123844 50764 123900
rect 50820 123844 50848 123900
rect 50528 122332 50848 123844
rect 50528 122276 50556 122332
rect 50612 122276 50660 122332
rect 50716 122276 50764 122332
rect 50820 122276 50848 122332
rect 50528 120764 50848 122276
rect 50528 120708 50556 120764
rect 50612 120708 50660 120764
rect 50716 120708 50764 120764
rect 50820 120708 50848 120764
rect 50528 119196 50848 120708
rect 50528 119140 50556 119196
rect 50612 119140 50660 119196
rect 50716 119140 50764 119196
rect 50820 119140 50848 119196
rect 50528 117628 50848 119140
rect 50528 117572 50556 117628
rect 50612 117572 50660 117628
rect 50716 117572 50764 117628
rect 50820 117572 50848 117628
rect 50528 116060 50848 117572
rect 50528 116004 50556 116060
rect 50612 116004 50660 116060
rect 50716 116004 50764 116060
rect 50820 116004 50848 116060
rect 50528 114492 50848 116004
rect 50528 114436 50556 114492
rect 50612 114436 50660 114492
rect 50716 114436 50764 114492
rect 50820 114436 50848 114492
rect 50528 112924 50848 114436
rect 50528 112868 50556 112924
rect 50612 112868 50660 112924
rect 50716 112868 50764 112924
rect 50820 112868 50848 112924
rect 50528 111356 50848 112868
rect 50528 111300 50556 111356
rect 50612 111300 50660 111356
rect 50716 111300 50764 111356
rect 50820 111300 50848 111356
rect 50528 109788 50848 111300
rect 50528 109732 50556 109788
rect 50612 109732 50660 109788
rect 50716 109732 50764 109788
rect 50820 109732 50848 109788
rect 50528 108220 50848 109732
rect 50528 108164 50556 108220
rect 50612 108164 50660 108220
rect 50716 108164 50764 108220
rect 50820 108164 50848 108220
rect 50528 106652 50848 108164
rect 50528 106596 50556 106652
rect 50612 106596 50660 106652
rect 50716 106596 50764 106652
rect 50820 106596 50848 106652
rect 50528 105084 50848 106596
rect 50528 105028 50556 105084
rect 50612 105028 50660 105084
rect 50716 105028 50764 105084
rect 50820 105028 50848 105084
rect 50528 103516 50848 105028
rect 50528 103460 50556 103516
rect 50612 103460 50660 103516
rect 50716 103460 50764 103516
rect 50820 103460 50848 103516
rect 50528 101948 50848 103460
rect 50528 101892 50556 101948
rect 50612 101892 50660 101948
rect 50716 101892 50764 101948
rect 50820 101892 50848 101948
rect 50528 100380 50848 101892
rect 50528 100324 50556 100380
rect 50612 100324 50660 100380
rect 50716 100324 50764 100380
rect 50820 100324 50848 100380
rect 50528 98812 50848 100324
rect 50528 98756 50556 98812
rect 50612 98756 50660 98812
rect 50716 98756 50764 98812
rect 50820 98756 50848 98812
rect 50528 97244 50848 98756
rect 50528 97188 50556 97244
rect 50612 97188 50660 97244
rect 50716 97188 50764 97244
rect 50820 97188 50848 97244
rect 50528 95676 50848 97188
rect 50528 95620 50556 95676
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50820 95620 50848 95676
rect 50528 94108 50848 95620
rect 50528 94052 50556 94108
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50820 94052 50848 94108
rect 50528 92540 50848 94052
rect 50528 92484 50556 92540
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50820 92484 50848 92540
rect 50528 90972 50848 92484
rect 50528 90916 50556 90972
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50820 90916 50848 90972
rect 50528 89404 50848 90916
rect 50528 89348 50556 89404
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50820 89348 50848 89404
rect 50528 87836 50848 89348
rect 50528 87780 50556 87836
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50820 87780 50848 87836
rect 50528 86268 50848 87780
rect 50528 86212 50556 86268
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50820 86212 50848 86268
rect 50528 84700 50848 86212
rect 50528 84644 50556 84700
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50820 84644 50848 84700
rect 50528 83132 50848 84644
rect 50528 83076 50556 83132
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50820 83076 50848 83132
rect 50528 81564 50848 83076
rect 50528 81508 50556 81564
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50820 81508 50848 81564
rect 50528 79996 50848 81508
rect 50528 79940 50556 79996
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50820 79940 50848 79996
rect 50528 78428 50848 79940
rect 50528 78372 50556 78428
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50820 78372 50848 78428
rect 50528 76860 50848 78372
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 132524 66208 132556
rect 65888 132468 65916 132524
rect 65972 132468 66020 132524
rect 66076 132468 66124 132524
rect 66180 132468 66208 132524
rect 65888 130956 66208 132468
rect 65888 130900 65916 130956
rect 65972 130900 66020 130956
rect 66076 130900 66124 130956
rect 66180 130900 66208 130956
rect 65888 129388 66208 130900
rect 65888 129332 65916 129388
rect 65972 129332 66020 129388
rect 66076 129332 66124 129388
rect 66180 129332 66208 129388
rect 65888 127820 66208 129332
rect 65888 127764 65916 127820
rect 65972 127764 66020 127820
rect 66076 127764 66124 127820
rect 66180 127764 66208 127820
rect 65888 126252 66208 127764
rect 65888 126196 65916 126252
rect 65972 126196 66020 126252
rect 66076 126196 66124 126252
rect 66180 126196 66208 126252
rect 65888 124684 66208 126196
rect 65888 124628 65916 124684
rect 65972 124628 66020 124684
rect 66076 124628 66124 124684
rect 66180 124628 66208 124684
rect 65888 123116 66208 124628
rect 65888 123060 65916 123116
rect 65972 123060 66020 123116
rect 66076 123060 66124 123116
rect 66180 123060 66208 123116
rect 65888 121548 66208 123060
rect 65888 121492 65916 121548
rect 65972 121492 66020 121548
rect 66076 121492 66124 121548
rect 66180 121492 66208 121548
rect 65888 119980 66208 121492
rect 65888 119924 65916 119980
rect 65972 119924 66020 119980
rect 66076 119924 66124 119980
rect 66180 119924 66208 119980
rect 65888 118412 66208 119924
rect 65888 118356 65916 118412
rect 65972 118356 66020 118412
rect 66076 118356 66124 118412
rect 66180 118356 66208 118412
rect 65888 116844 66208 118356
rect 65888 116788 65916 116844
rect 65972 116788 66020 116844
rect 66076 116788 66124 116844
rect 66180 116788 66208 116844
rect 65888 115276 66208 116788
rect 65888 115220 65916 115276
rect 65972 115220 66020 115276
rect 66076 115220 66124 115276
rect 66180 115220 66208 115276
rect 65888 113708 66208 115220
rect 65888 113652 65916 113708
rect 65972 113652 66020 113708
rect 66076 113652 66124 113708
rect 66180 113652 66208 113708
rect 65888 112140 66208 113652
rect 65888 112084 65916 112140
rect 65972 112084 66020 112140
rect 66076 112084 66124 112140
rect 66180 112084 66208 112140
rect 65888 110572 66208 112084
rect 65888 110516 65916 110572
rect 65972 110516 66020 110572
rect 66076 110516 66124 110572
rect 66180 110516 66208 110572
rect 65888 109004 66208 110516
rect 65888 108948 65916 109004
rect 65972 108948 66020 109004
rect 66076 108948 66124 109004
rect 66180 108948 66208 109004
rect 65888 107436 66208 108948
rect 65888 107380 65916 107436
rect 65972 107380 66020 107436
rect 66076 107380 66124 107436
rect 66180 107380 66208 107436
rect 65888 105868 66208 107380
rect 65888 105812 65916 105868
rect 65972 105812 66020 105868
rect 66076 105812 66124 105868
rect 66180 105812 66208 105868
rect 65888 104300 66208 105812
rect 65888 104244 65916 104300
rect 65972 104244 66020 104300
rect 66076 104244 66124 104300
rect 66180 104244 66208 104300
rect 65888 102732 66208 104244
rect 65888 102676 65916 102732
rect 65972 102676 66020 102732
rect 66076 102676 66124 102732
rect 66180 102676 66208 102732
rect 65888 101164 66208 102676
rect 65888 101108 65916 101164
rect 65972 101108 66020 101164
rect 66076 101108 66124 101164
rect 66180 101108 66208 101164
rect 65888 99596 66208 101108
rect 65888 99540 65916 99596
rect 65972 99540 66020 99596
rect 66076 99540 66124 99596
rect 66180 99540 66208 99596
rect 65888 98028 66208 99540
rect 65888 97972 65916 98028
rect 65972 97972 66020 98028
rect 66076 97972 66124 98028
rect 66180 97972 66208 98028
rect 65888 96460 66208 97972
rect 65888 96404 65916 96460
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 66180 96404 66208 96460
rect 65888 94892 66208 96404
rect 65888 94836 65916 94892
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 66180 94836 66208 94892
rect 65888 93324 66208 94836
rect 65888 93268 65916 93324
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 66180 93268 66208 93324
rect 65888 91756 66208 93268
rect 65888 91700 65916 91756
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 66180 91700 66208 91756
rect 65888 90188 66208 91700
rect 65888 90132 65916 90188
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 66180 90132 66208 90188
rect 65888 88620 66208 90132
rect 65888 88564 65916 88620
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 66180 88564 66208 88620
rect 65888 87052 66208 88564
rect 65888 86996 65916 87052
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 66180 86996 66208 87052
rect 65888 85484 66208 86996
rect 65888 85428 65916 85484
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 66180 85428 66208 85484
rect 65888 83916 66208 85428
rect 65888 83860 65916 83916
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 66180 83860 66208 83916
rect 65888 82348 66208 83860
rect 65888 82292 65916 82348
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 66180 82292 66208 82348
rect 65888 80780 66208 82292
rect 65888 80724 65916 80780
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 66180 80724 66208 80780
rect 65888 79212 66208 80724
rect 65888 79156 65916 79212
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 66180 79156 66208 79212
rect 65888 77644 66208 79156
rect 65888 77588 65916 77644
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 66180 77588 66208 77644
rect 65888 76076 66208 77588
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
rect 81248 131740 81568 132556
rect 81248 131684 81276 131740
rect 81332 131684 81380 131740
rect 81436 131684 81484 131740
rect 81540 131684 81568 131740
rect 81248 130172 81568 131684
rect 81248 130116 81276 130172
rect 81332 130116 81380 130172
rect 81436 130116 81484 130172
rect 81540 130116 81568 130172
rect 81248 128604 81568 130116
rect 81248 128548 81276 128604
rect 81332 128548 81380 128604
rect 81436 128548 81484 128604
rect 81540 128548 81568 128604
rect 81248 127036 81568 128548
rect 81248 126980 81276 127036
rect 81332 126980 81380 127036
rect 81436 126980 81484 127036
rect 81540 126980 81568 127036
rect 81248 125468 81568 126980
rect 81248 125412 81276 125468
rect 81332 125412 81380 125468
rect 81436 125412 81484 125468
rect 81540 125412 81568 125468
rect 81248 123900 81568 125412
rect 81248 123844 81276 123900
rect 81332 123844 81380 123900
rect 81436 123844 81484 123900
rect 81540 123844 81568 123900
rect 81248 122332 81568 123844
rect 81248 122276 81276 122332
rect 81332 122276 81380 122332
rect 81436 122276 81484 122332
rect 81540 122276 81568 122332
rect 81248 120764 81568 122276
rect 81248 120708 81276 120764
rect 81332 120708 81380 120764
rect 81436 120708 81484 120764
rect 81540 120708 81568 120764
rect 81248 119196 81568 120708
rect 81248 119140 81276 119196
rect 81332 119140 81380 119196
rect 81436 119140 81484 119196
rect 81540 119140 81568 119196
rect 81248 117628 81568 119140
rect 81248 117572 81276 117628
rect 81332 117572 81380 117628
rect 81436 117572 81484 117628
rect 81540 117572 81568 117628
rect 81248 116060 81568 117572
rect 81248 116004 81276 116060
rect 81332 116004 81380 116060
rect 81436 116004 81484 116060
rect 81540 116004 81568 116060
rect 81248 114492 81568 116004
rect 81248 114436 81276 114492
rect 81332 114436 81380 114492
rect 81436 114436 81484 114492
rect 81540 114436 81568 114492
rect 81248 112924 81568 114436
rect 81248 112868 81276 112924
rect 81332 112868 81380 112924
rect 81436 112868 81484 112924
rect 81540 112868 81568 112924
rect 81248 111356 81568 112868
rect 81248 111300 81276 111356
rect 81332 111300 81380 111356
rect 81436 111300 81484 111356
rect 81540 111300 81568 111356
rect 81248 109788 81568 111300
rect 81248 109732 81276 109788
rect 81332 109732 81380 109788
rect 81436 109732 81484 109788
rect 81540 109732 81568 109788
rect 81248 108220 81568 109732
rect 81248 108164 81276 108220
rect 81332 108164 81380 108220
rect 81436 108164 81484 108220
rect 81540 108164 81568 108220
rect 81248 106652 81568 108164
rect 81248 106596 81276 106652
rect 81332 106596 81380 106652
rect 81436 106596 81484 106652
rect 81540 106596 81568 106652
rect 81248 105084 81568 106596
rect 81248 105028 81276 105084
rect 81332 105028 81380 105084
rect 81436 105028 81484 105084
rect 81540 105028 81568 105084
rect 81248 103516 81568 105028
rect 81248 103460 81276 103516
rect 81332 103460 81380 103516
rect 81436 103460 81484 103516
rect 81540 103460 81568 103516
rect 81248 101948 81568 103460
rect 81248 101892 81276 101948
rect 81332 101892 81380 101948
rect 81436 101892 81484 101948
rect 81540 101892 81568 101948
rect 81248 100380 81568 101892
rect 81248 100324 81276 100380
rect 81332 100324 81380 100380
rect 81436 100324 81484 100380
rect 81540 100324 81568 100380
rect 81248 98812 81568 100324
rect 81248 98756 81276 98812
rect 81332 98756 81380 98812
rect 81436 98756 81484 98812
rect 81540 98756 81568 98812
rect 81248 97244 81568 98756
rect 81248 97188 81276 97244
rect 81332 97188 81380 97244
rect 81436 97188 81484 97244
rect 81540 97188 81568 97244
rect 81248 95676 81568 97188
rect 81248 95620 81276 95676
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81540 95620 81568 95676
rect 81248 94108 81568 95620
rect 81248 94052 81276 94108
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81540 94052 81568 94108
rect 81248 92540 81568 94052
rect 81248 92484 81276 92540
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81540 92484 81568 92540
rect 81248 90972 81568 92484
rect 81248 90916 81276 90972
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81540 90916 81568 90972
rect 81248 89404 81568 90916
rect 81248 89348 81276 89404
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81540 89348 81568 89404
rect 81248 87836 81568 89348
rect 81248 87780 81276 87836
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81540 87780 81568 87836
rect 81248 86268 81568 87780
rect 81248 86212 81276 86268
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81540 86212 81568 86268
rect 81248 84700 81568 86212
rect 81248 84644 81276 84700
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81540 84644 81568 84700
rect 81248 83132 81568 84644
rect 81248 83076 81276 83132
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81540 83076 81568 83132
rect 81248 81564 81568 83076
rect 81248 81508 81276 81564
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81540 81508 81568 81564
rect 81248 79996 81568 81508
rect 81248 79940 81276 79996
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81540 79940 81568 79996
rect 81248 78428 81568 79940
rect 81248 78372 81276 78428
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81540 78372 81568 78428
rect 81248 76860 81568 78372
rect 81248 76804 81276 76860
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81540 76804 81568 76860
rect 81248 75292 81568 76804
rect 81248 75236 81276 75292
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81540 75236 81568 75292
rect 81248 73724 81568 75236
rect 81248 73668 81276 73724
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81540 73668 81568 73724
rect 81248 72156 81568 73668
rect 81248 72100 81276 72156
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81540 72100 81568 72156
rect 81248 70588 81568 72100
rect 81248 70532 81276 70588
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81540 70532 81568 70588
rect 81248 69020 81568 70532
rect 81248 68964 81276 69020
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81540 68964 81568 69020
rect 81248 67452 81568 68964
rect 81248 67396 81276 67452
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81540 67396 81568 67452
rect 81248 65884 81568 67396
rect 81248 65828 81276 65884
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81540 65828 81568 65884
rect 81248 64316 81568 65828
rect 81248 64260 81276 64316
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81540 64260 81568 64316
rect 81248 62748 81568 64260
rect 81248 62692 81276 62748
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81540 62692 81568 62748
rect 81248 61180 81568 62692
rect 81248 61124 81276 61180
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81540 61124 81568 61180
rect 81248 59612 81568 61124
rect 81248 59556 81276 59612
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81540 59556 81568 59612
rect 81248 58044 81568 59556
rect 81248 57988 81276 58044
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81540 57988 81568 58044
rect 81248 56476 81568 57988
rect 81248 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81568 56476
rect 81248 54908 81568 56420
rect 81248 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81568 54908
rect 81248 53340 81568 54852
rect 81248 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81568 53340
rect 81248 51772 81568 53284
rect 81248 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81568 51772
rect 81248 50204 81568 51716
rect 81248 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81568 50204
rect 81248 48636 81568 50148
rect 81248 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81568 48636
rect 81248 47068 81568 48580
rect 81248 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81568 47068
rect 81248 45500 81568 47012
rect 81248 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81568 45500
rect 81248 43932 81568 45444
rect 81248 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81568 43932
rect 81248 42364 81568 43876
rect 81248 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81568 42364
rect 81248 40796 81568 42308
rect 81248 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81568 40796
rect 81248 39228 81568 40740
rect 81248 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81568 39228
rect 81248 37660 81568 39172
rect 81248 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81568 37660
rect 81248 36092 81568 37604
rect 81248 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81568 36092
rect 81248 34524 81568 36036
rect 81248 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81568 34524
rect 81248 32956 81568 34468
rect 81248 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81568 32956
rect 81248 31388 81568 32900
rect 81248 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81568 31388
rect 81248 29820 81568 31332
rect 81248 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81568 29820
rect 81248 28252 81568 29764
rect 81248 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81568 28252
rect 81248 26684 81568 28196
rect 81248 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81568 26684
rect 81248 25116 81568 26628
rect 81248 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81568 25116
rect 81248 23548 81568 25060
rect 81248 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81568 23548
rect 81248 21980 81568 23492
rect 81248 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81568 21980
rect 81248 20412 81568 21924
rect 81248 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81568 20412
rect 81248 18844 81568 20356
rect 81248 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81568 18844
rect 81248 17276 81568 18788
rect 81248 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81568 17276
rect 81248 15708 81568 17220
rect 81248 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81568 15708
rect 81248 14140 81568 15652
rect 81248 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81568 14140
rect 81248 12572 81568 14084
rect 81248 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81568 12572
rect 81248 11004 81568 12516
rect 81248 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81568 11004
rect 81248 9436 81568 10948
rect 81248 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81568 9436
rect 81248 7868 81568 9380
rect 81248 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81568 7868
rect 81248 6300 81568 7812
rect 81248 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81568 6300
rect 81248 4732 81568 6244
rect 81248 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81568 4732
rect 81248 3164 81568 4676
rect 81248 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81568 3164
rect 81248 3076 81568 3108
rect 96608 132524 96928 132556
rect 96608 132468 96636 132524
rect 96692 132468 96740 132524
rect 96796 132468 96844 132524
rect 96900 132468 96928 132524
rect 96608 130956 96928 132468
rect 96608 130900 96636 130956
rect 96692 130900 96740 130956
rect 96796 130900 96844 130956
rect 96900 130900 96928 130956
rect 96608 129388 96928 130900
rect 96608 129332 96636 129388
rect 96692 129332 96740 129388
rect 96796 129332 96844 129388
rect 96900 129332 96928 129388
rect 96608 127820 96928 129332
rect 96608 127764 96636 127820
rect 96692 127764 96740 127820
rect 96796 127764 96844 127820
rect 96900 127764 96928 127820
rect 96608 126252 96928 127764
rect 96608 126196 96636 126252
rect 96692 126196 96740 126252
rect 96796 126196 96844 126252
rect 96900 126196 96928 126252
rect 96608 124684 96928 126196
rect 96608 124628 96636 124684
rect 96692 124628 96740 124684
rect 96796 124628 96844 124684
rect 96900 124628 96928 124684
rect 96608 123116 96928 124628
rect 96608 123060 96636 123116
rect 96692 123060 96740 123116
rect 96796 123060 96844 123116
rect 96900 123060 96928 123116
rect 96608 121548 96928 123060
rect 96608 121492 96636 121548
rect 96692 121492 96740 121548
rect 96796 121492 96844 121548
rect 96900 121492 96928 121548
rect 96608 119980 96928 121492
rect 96608 119924 96636 119980
rect 96692 119924 96740 119980
rect 96796 119924 96844 119980
rect 96900 119924 96928 119980
rect 96608 118412 96928 119924
rect 96608 118356 96636 118412
rect 96692 118356 96740 118412
rect 96796 118356 96844 118412
rect 96900 118356 96928 118412
rect 96608 116844 96928 118356
rect 96608 116788 96636 116844
rect 96692 116788 96740 116844
rect 96796 116788 96844 116844
rect 96900 116788 96928 116844
rect 96608 115276 96928 116788
rect 96608 115220 96636 115276
rect 96692 115220 96740 115276
rect 96796 115220 96844 115276
rect 96900 115220 96928 115276
rect 96608 113708 96928 115220
rect 96608 113652 96636 113708
rect 96692 113652 96740 113708
rect 96796 113652 96844 113708
rect 96900 113652 96928 113708
rect 96608 112140 96928 113652
rect 96608 112084 96636 112140
rect 96692 112084 96740 112140
rect 96796 112084 96844 112140
rect 96900 112084 96928 112140
rect 96608 110572 96928 112084
rect 96608 110516 96636 110572
rect 96692 110516 96740 110572
rect 96796 110516 96844 110572
rect 96900 110516 96928 110572
rect 96608 109004 96928 110516
rect 96608 108948 96636 109004
rect 96692 108948 96740 109004
rect 96796 108948 96844 109004
rect 96900 108948 96928 109004
rect 96608 107436 96928 108948
rect 96608 107380 96636 107436
rect 96692 107380 96740 107436
rect 96796 107380 96844 107436
rect 96900 107380 96928 107436
rect 96608 105868 96928 107380
rect 96608 105812 96636 105868
rect 96692 105812 96740 105868
rect 96796 105812 96844 105868
rect 96900 105812 96928 105868
rect 96608 104300 96928 105812
rect 96608 104244 96636 104300
rect 96692 104244 96740 104300
rect 96796 104244 96844 104300
rect 96900 104244 96928 104300
rect 96608 102732 96928 104244
rect 96608 102676 96636 102732
rect 96692 102676 96740 102732
rect 96796 102676 96844 102732
rect 96900 102676 96928 102732
rect 96608 101164 96928 102676
rect 96608 101108 96636 101164
rect 96692 101108 96740 101164
rect 96796 101108 96844 101164
rect 96900 101108 96928 101164
rect 96608 99596 96928 101108
rect 96608 99540 96636 99596
rect 96692 99540 96740 99596
rect 96796 99540 96844 99596
rect 96900 99540 96928 99596
rect 96608 98028 96928 99540
rect 96608 97972 96636 98028
rect 96692 97972 96740 98028
rect 96796 97972 96844 98028
rect 96900 97972 96928 98028
rect 96608 96460 96928 97972
rect 96608 96404 96636 96460
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96900 96404 96928 96460
rect 96608 94892 96928 96404
rect 96608 94836 96636 94892
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96900 94836 96928 94892
rect 96608 93324 96928 94836
rect 96608 93268 96636 93324
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96900 93268 96928 93324
rect 96608 91756 96928 93268
rect 96608 91700 96636 91756
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96900 91700 96928 91756
rect 96608 90188 96928 91700
rect 96608 90132 96636 90188
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96900 90132 96928 90188
rect 96608 88620 96928 90132
rect 96608 88564 96636 88620
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96900 88564 96928 88620
rect 96608 87052 96928 88564
rect 96608 86996 96636 87052
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96900 86996 96928 87052
rect 96608 85484 96928 86996
rect 96608 85428 96636 85484
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96900 85428 96928 85484
rect 96608 83916 96928 85428
rect 96608 83860 96636 83916
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96900 83860 96928 83916
rect 96608 82348 96928 83860
rect 96608 82292 96636 82348
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96900 82292 96928 82348
rect 96608 80780 96928 82292
rect 96608 80724 96636 80780
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96900 80724 96928 80780
rect 96608 79212 96928 80724
rect 96608 79156 96636 79212
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96900 79156 96928 79212
rect 96608 77644 96928 79156
rect 96608 77588 96636 77644
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96900 77588 96928 77644
rect 96608 76076 96928 77588
rect 96608 76020 96636 76076
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96900 76020 96928 76076
rect 96608 74508 96928 76020
rect 96608 74452 96636 74508
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96900 74452 96928 74508
rect 96608 72940 96928 74452
rect 96608 72884 96636 72940
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96900 72884 96928 72940
rect 96608 71372 96928 72884
rect 96608 71316 96636 71372
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96900 71316 96928 71372
rect 96608 69804 96928 71316
rect 96608 69748 96636 69804
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96900 69748 96928 69804
rect 96608 68236 96928 69748
rect 96608 68180 96636 68236
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96900 68180 96928 68236
rect 96608 66668 96928 68180
rect 96608 66612 96636 66668
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96900 66612 96928 66668
rect 96608 65100 96928 66612
rect 96608 65044 96636 65100
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96900 65044 96928 65100
rect 96608 63532 96928 65044
rect 96608 63476 96636 63532
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96900 63476 96928 63532
rect 96608 61964 96928 63476
rect 96608 61908 96636 61964
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96900 61908 96928 61964
rect 96608 60396 96928 61908
rect 96608 60340 96636 60396
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96900 60340 96928 60396
rect 96608 58828 96928 60340
rect 96608 58772 96636 58828
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96900 58772 96928 58828
rect 96608 57260 96928 58772
rect 96608 57204 96636 57260
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96900 57204 96928 57260
rect 96608 55692 96928 57204
rect 96608 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96928 55692
rect 96608 54124 96928 55636
rect 96608 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96928 54124
rect 96608 52556 96928 54068
rect 96608 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96928 52556
rect 96608 50988 96928 52500
rect 96608 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96928 50988
rect 96608 49420 96928 50932
rect 96608 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96928 49420
rect 96608 47852 96928 49364
rect 96608 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96928 47852
rect 96608 46284 96928 47796
rect 96608 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96928 46284
rect 96608 44716 96928 46228
rect 96608 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96928 44716
rect 96608 43148 96928 44660
rect 96608 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96928 43148
rect 96608 41580 96928 43092
rect 96608 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96928 41580
rect 96608 40012 96928 41524
rect 96608 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96928 40012
rect 96608 38444 96928 39956
rect 96608 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96928 38444
rect 96608 36876 96928 38388
rect 96608 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96928 36876
rect 96608 35308 96928 36820
rect 96608 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96928 35308
rect 96608 33740 96928 35252
rect 96608 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96928 33740
rect 96608 32172 96928 33684
rect 96608 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96928 32172
rect 96608 30604 96928 32116
rect 96608 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96928 30604
rect 96608 29036 96928 30548
rect 96608 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96928 29036
rect 96608 27468 96928 28980
rect 96608 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96928 27468
rect 96608 25900 96928 27412
rect 96608 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96928 25900
rect 96608 24332 96928 25844
rect 96608 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96928 24332
rect 96608 22764 96928 24276
rect 96608 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96928 22764
rect 96608 21196 96928 22708
rect 96608 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96928 21196
rect 96608 19628 96928 21140
rect 96608 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96928 19628
rect 96608 18060 96928 19572
rect 96608 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96928 18060
rect 96608 16492 96928 18004
rect 96608 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96928 16492
rect 96608 14924 96928 16436
rect 96608 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96928 14924
rect 96608 13356 96928 14868
rect 96608 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96928 13356
rect 96608 11788 96928 13300
rect 96608 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96928 11788
rect 96608 10220 96928 11732
rect 96608 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96928 10220
rect 96608 8652 96928 10164
rect 96608 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96928 8652
rect 96608 7084 96928 8596
rect 96608 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96928 7084
rect 96608 5516 96928 7028
rect 96608 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96928 5516
rect 96608 3948 96928 5460
rect 96608 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96928 3948
rect 96608 3076 96928 3892
rect 111968 131740 112288 132556
rect 111968 131684 111996 131740
rect 112052 131684 112100 131740
rect 112156 131684 112204 131740
rect 112260 131684 112288 131740
rect 111968 130172 112288 131684
rect 111968 130116 111996 130172
rect 112052 130116 112100 130172
rect 112156 130116 112204 130172
rect 112260 130116 112288 130172
rect 111968 128604 112288 130116
rect 111968 128548 111996 128604
rect 112052 128548 112100 128604
rect 112156 128548 112204 128604
rect 112260 128548 112288 128604
rect 111968 127036 112288 128548
rect 111968 126980 111996 127036
rect 112052 126980 112100 127036
rect 112156 126980 112204 127036
rect 112260 126980 112288 127036
rect 111968 125468 112288 126980
rect 111968 125412 111996 125468
rect 112052 125412 112100 125468
rect 112156 125412 112204 125468
rect 112260 125412 112288 125468
rect 111968 123900 112288 125412
rect 111968 123844 111996 123900
rect 112052 123844 112100 123900
rect 112156 123844 112204 123900
rect 112260 123844 112288 123900
rect 111968 122332 112288 123844
rect 111968 122276 111996 122332
rect 112052 122276 112100 122332
rect 112156 122276 112204 122332
rect 112260 122276 112288 122332
rect 111968 120764 112288 122276
rect 111968 120708 111996 120764
rect 112052 120708 112100 120764
rect 112156 120708 112204 120764
rect 112260 120708 112288 120764
rect 111968 119196 112288 120708
rect 111968 119140 111996 119196
rect 112052 119140 112100 119196
rect 112156 119140 112204 119196
rect 112260 119140 112288 119196
rect 111968 117628 112288 119140
rect 111968 117572 111996 117628
rect 112052 117572 112100 117628
rect 112156 117572 112204 117628
rect 112260 117572 112288 117628
rect 111968 116060 112288 117572
rect 111968 116004 111996 116060
rect 112052 116004 112100 116060
rect 112156 116004 112204 116060
rect 112260 116004 112288 116060
rect 111968 114492 112288 116004
rect 111968 114436 111996 114492
rect 112052 114436 112100 114492
rect 112156 114436 112204 114492
rect 112260 114436 112288 114492
rect 111968 112924 112288 114436
rect 111968 112868 111996 112924
rect 112052 112868 112100 112924
rect 112156 112868 112204 112924
rect 112260 112868 112288 112924
rect 111968 111356 112288 112868
rect 111968 111300 111996 111356
rect 112052 111300 112100 111356
rect 112156 111300 112204 111356
rect 112260 111300 112288 111356
rect 111968 109788 112288 111300
rect 111968 109732 111996 109788
rect 112052 109732 112100 109788
rect 112156 109732 112204 109788
rect 112260 109732 112288 109788
rect 111968 108220 112288 109732
rect 111968 108164 111996 108220
rect 112052 108164 112100 108220
rect 112156 108164 112204 108220
rect 112260 108164 112288 108220
rect 111968 106652 112288 108164
rect 111968 106596 111996 106652
rect 112052 106596 112100 106652
rect 112156 106596 112204 106652
rect 112260 106596 112288 106652
rect 111968 105084 112288 106596
rect 111968 105028 111996 105084
rect 112052 105028 112100 105084
rect 112156 105028 112204 105084
rect 112260 105028 112288 105084
rect 111968 103516 112288 105028
rect 111968 103460 111996 103516
rect 112052 103460 112100 103516
rect 112156 103460 112204 103516
rect 112260 103460 112288 103516
rect 111968 101948 112288 103460
rect 111968 101892 111996 101948
rect 112052 101892 112100 101948
rect 112156 101892 112204 101948
rect 112260 101892 112288 101948
rect 111968 100380 112288 101892
rect 111968 100324 111996 100380
rect 112052 100324 112100 100380
rect 112156 100324 112204 100380
rect 112260 100324 112288 100380
rect 111968 98812 112288 100324
rect 111968 98756 111996 98812
rect 112052 98756 112100 98812
rect 112156 98756 112204 98812
rect 112260 98756 112288 98812
rect 111968 97244 112288 98756
rect 111968 97188 111996 97244
rect 112052 97188 112100 97244
rect 112156 97188 112204 97244
rect 112260 97188 112288 97244
rect 111968 95676 112288 97188
rect 111968 95620 111996 95676
rect 112052 95620 112100 95676
rect 112156 95620 112204 95676
rect 112260 95620 112288 95676
rect 111968 94108 112288 95620
rect 111968 94052 111996 94108
rect 112052 94052 112100 94108
rect 112156 94052 112204 94108
rect 112260 94052 112288 94108
rect 111968 92540 112288 94052
rect 111968 92484 111996 92540
rect 112052 92484 112100 92540
rect 112156 92484 112204 92540
rect 112260 92484 112288 92540
rect 111968 90972 112288 92484
rect 111968 90916 111996 90972
rect 112052 90916 112100 90972
rect 112156 90916 112204 90972
rect 112260 90916 112288 90972
rect 111968 89404 112288 90916
rect 111968 89348 111996 89404
rect 112052 89348 112100 89404
rect 112156 89348 112204 89404
rect 112260 89348 112288 89404
rect 111968 87836 112288 89348
rect 111968 87780 111996 87836
rect 112052 87780 112100 87836
rect 112156 87780 112204 87836
rect 112260 87780 112288 87836
rect 111968 86268 112288 87780
rect 111968 86212 111996 86268
rect 112052 86212 112100 86268
rect 112156 86212 112204 86268
rect 112260 86212 112288 86268
rect 111968 84700 112288 86212
rect 111968 84644 111996 84700
rect 112052 84644 112100 84700
rect 112156 84644 112204 84700
rect 112260 84644 112288 84700
rect 111968 83132 112288 84644
rect 111968 83076 111996 83132
rect 112052 83076 112100 83132
rect 112156 83076 112204 83132
rect 112260 83076 112288 83132
rect 111968 81564 112288 83076
rect 111968 81508 111996 81564
rect 112052 81508 112100 81564
rect 112156 81508 112204 81564
rect 112260 81508 112288 81564
rect 111968 79996 112288 81508
rect 111968 79940 111996 79996
rect 112052 79940 112100 79996
rect 112156 79940 112204 79996
rect 112260 79940 112288 79996
rect 111968 78428 112288 79940
rect 111968 78372 111996 78428
rect 112052 78372 112100 78428
rect 112156 78372 112204 78428
rect 112260 78372 112288 78428
rect 111968 76860 112288 78372
rect 111968 76804 111996 76860
rect 112052 76804 112100 76860
rect 112156 76804 112204 76860
rect 112260 76804 112288 76860
rect 111968 75292 112288 76804
rect 111968 75236 111996 75292
rect 112052 75236 112100 75292
rect 112156 75236 112204 75292
rect 112260 75236 112288 75292
rect 111968 73724 112288 75236
rect 111968 73668 111996 73724
rect 112052 73668 112100 73724
rect 112156 73668 112204 73724
rect 112260 73668 112288 73724
rect 111968 72156 112288 73668
rect 111968 72100 111996 72156
rect 112052 72100 112100 72156
rect 112156 72100 112204 72156
rect 112260 72100 112288 72156
rect 111968 70588 112288 72100
rect 111968 70532 111996 70588
rect 112052 70532 112100 70588
rect 112156 70532 112204 70588
rect 112260 70532 112288 70588
rect 111968 69020 112288 70532
rect 111968 68964 111996 69020
rect 112052 68964 112100 69020
rect 112156 68964 112204 69020
rect 112260 68964 112288 69020
rect 111968 67452 112288 68964
rect 111968 67396 111996 67452
rect 112052 67396 112100 67452
rect 112156 67396 112204 67452
rect 112260 67396 112288 67452
rect 111968 65884 112288 67396
rect 111968 65828 111996 65884
rect 112052 65828 112100 65884
rect 112156 65828 112204 65884
rect 112260 65828 112288 65884
rect 111968 64316 112288 65828
rect 111968 64260 111996 64316
rect 112052 64260 112100 64316
rect 112156 64260 112204 64316
rect 112260 64260 112288 64316
rect 111968 62748 112288 64260
rect 111968 62692 111996 62748
rect 112052 62692 112100 62748
rect 112156 62692 112204 62748
rect 112260 62692 112288 62748
rect 111968 61180 112288 62692
rect 111968 61124 111996 61180
rect 112052 61124 112100 61180
rect 112156 61124 112204 61180
rect 112260 61124 112288 61180
rect 111968 59612 112288 61124
rect 111968 59556 111996 59612
rect 112052 59556 112100 59612
rect 112156 59556 112204 59612
rect 112260 59556 112288 59612
rect 111968 58044 112288 59556
rect 111968 57988 111996 58044
rect 112052 57988 112100 58044
rect 112156 57988 112204 58044
rect 112260 57988 112288 58044
rect 111968 56476 112288 57988
rect 111968 56420 111996 56476
rect 112052 56420 112100 56476
rect 112156 56420 112204 56476
rect 112260 56420 112288 56476
rect 111968 54908 112288 56420
rect 111968 54852 111996 54908
rect 112052 54852 112100 54908
rect 112156 54852 112204 54908
rect 112260 54852 112288 54908
rect 111968 53340 112288 54852
rect 111968 53284 111996 53340
rect 112052 53284 112100 53340
rect 112156 53284 112204 53340
rect 112260 53284 112288 53340
rect 111968 51772 112288 53284
rect 111968 51716 111996 51772
rect 112052 51716 112100 51772
rect 112156 51716 112204 51772
rect 112260 51716 112288 51772
rect 111968 50204 112288 51716
rect 111968 50148 111996 50204
rect 112052 50148 112100 50204
rect 112156 50148 112204 50204
rect 112260 50148 112288 50204
rect 111968 48636 112288 50148
rect 111968 48580 111996 48636
rect 112052 48580 112100 48636
rect 112156 48580 112204 48636
rect 112260 48580 112288 48636
rect 111968 47068 112288 48580
rect 111968 47012 111996 47068
rect 112052 47012 112100 47068
rect 112156 47012 112204 47068
rect 112260 47012 112288 47068
rect 111968 45500 112288 47012
rect 111968 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112288 45500
rect 111968 43932 112288 45444
rect 111968 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112288 43932
rect 111968 42364 112288 43876
rect 111968 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112288 42364
rect 111968 40796 112288 42308
rect 111968 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112288 40796
rect 111968 39228 112288 40740
rect 111968 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112288 39228
rect 111968 37660 112288 39172
rect 111968 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112288 37660
rect 111968 36092 112288 37604
rect 111968 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112288 36092
rect 111968 34524 112288 36036
rect 111968 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112288 34524
rect 111968 32956 112288 34468
rect 111968 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112288 32956
rect 111968 31388 112288 32900
rect 111968 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112288 31388
rect 111968 29820 112288 31332
rect 111968 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112288 29820
rect 111968 28252 112288 29764
rect 111968 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112288 28252
rect 111968 26684 112288 28196
rect 111968 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112288 26684
rect 111968 25116 112288 26628
rect 111968 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112288 25116
rect 111968 23548 112288 25060
rect 111968 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112288 23548
rect 111968 21980 112288 23492
rect 111968 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112288 21980
rect 111968 20412 112288 21924
rect 111968 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112288 20412
rect 111968 18844 112288 20356
rect 111968 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112288 18844
rect 111968 17276 112288 18788
rect 111968 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112288 17276
rect 111968 15708 112288 17220
rect 111968 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112288 15708
rect 111968 14140 112288 15652
rect 111968 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112288 14140
rect 111968 12572 112288 14084
rect 111968 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112288 12572
rect 111968 11004 112288 12516
rect 111968 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112288 11004
rect 111968 9436 112288 10948
rect 111968 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112288 9436
rect 111968 7868 112288 9380
rect 111968 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112288 7868
rect 111968 6300 112288 7812
rect 111968 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112288 6300
rect 111968 4732 112288 6244
rect 111968 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112288 4732
rect 111968 3164 112288 4676
rect 111968 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112288 3164
rect 111968 3076 112288 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__002__I pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 3136 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__003__I
timestamp 1663859327
transform -1 0 20720 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__004__A2
timestamp 1663859327
transform 1 0 4032 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__005__CLK
timestamp 1663859327
transform 1 0 6272 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1663859327
transform -1 0 2128 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__I
timestamp 1663859327
transform 1 0 59360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I
timestamp 1663859327
transform 1 0 60032 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1663859327
transform -1 0 1904 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1663859327
transform -1 0 1904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1663859327
transform -1 0 1904 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1663859327
transform -1 0 1904 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1663859327
transform 1 0 2576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1663859327
transform 1 0 59808 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1663859327
transform -1 0 1904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output8_I
timestamp 1663859327
transform 1 0 116480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output9_I
timestamp 1663859327
transform 1 0 20608 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output10_I
timestamp 1663859327
transform 1 0 3472 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output11_I
timestamp 1663859327
transform 1 0 116256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output12_I
timestamp 1663859327
transform 1 0 3472 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2016 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2576 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 4368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37
timestamp 1663859327
transform 1 0 5488 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 7280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59
timestamp 1663859327
transform 1 0 7952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65
timestamp 1663859327
transform 1 0 8624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1663859327
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1663859327
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77
timestamp 1663859327
transform 1 0 9968 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93
timestamp 1663859327
transform 1 0 11760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101
timestamp 1663859327
transform 1 0 12656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1663859327
transform 1 0 13328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115
timestamp 1663859327
transform 1 0 14224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119
timestamp 1663859327
transform 1 0 14672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_125
timestamp 1663859327
transform 1 0 15344 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133
timestamp 1663859327
transform 1 0 16240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137
timestamp 1663859327
transform 1 0 16688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1663859327
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 17248 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1663859327
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_177
timestamp 1663859327
transform 1 0 21168 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1663859327
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_212
timestamp 1663859327
transform 1 0 25088 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_228
timestamp 1663859327
transform 1 0 26880 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_233
timestamp 1663859327
transform 1 0 27440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_237
timestamp 1663859327
transform 1 0 27888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_239
timestamp 1663859327
transform 1 0 28112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1663859327
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_247
timestamp 1663859327
transform 1 0 29008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_251
timestamp 1663859327
transform 1 0 29456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_257
timestamp 1663859327
transform 1 0 30128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_263
timestamp 1663859327
transform 1 0 30800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1663859327
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1663859327
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_287
timestamp 1663859327
transform 1 0 33488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_299
timestamp 1663859327
transform 1 0 34832 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317
timestamp 1663859327
transform 1 0 36848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_323
timestamp 1663859327
transform 1 0 37520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_329
timestamp 1663859327
transform 1 0 38192 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_345
timestamp 1663859327
transform 1 0 39984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1663859327
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_352
timestamp 1663859327
transform 1 0 40768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_368
timestamp 1663859327
transform 1 0 42560 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_372
timestamp 1663859327
transform 1 0 43008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_377
timestamp 1663859327
transform 1 0 43568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_387
timestamp 1663859327
transform 1 0 44688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_395
timestamp 1663859327
transform 1 0 45584 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_411
timestamp 1663859327
transform 1 0 47376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1663859327
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_422
timestamp 1663859327
transform 1 0 48608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_426
timestamp 1663859327
transform 1 0 49056 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_431
timestamp 1663859327
transform 1 0 49616 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_447
timestamp 1663859327
transform 1 0 51408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_449
timestamp 1663859327
transform 1 0 51632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1663859327
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1663859327
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_462
timestamp 1663859327
transform 1 0 53088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_466
timestamp 1663859327
transform 1 0 53536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_468
timestamp 1663859327
transform 1 0 53760 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_473
timestamp 1663859327
transform 1 0 54320 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_485
timestamp 1663859327
transform 1 0 55664 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1663859327
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_492
timestamp 1663859327
transform 1 0 56448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_508
timestamp 1663859327
transform 1 0 58240 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_516
timestamp 1663859327
transform 1 0 59136 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_521
timestamp 1663859327
transform 1 0 59696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_527
timestamp 1663859327
transform 1 0 60368 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_543
timestamp 1663859327
transform 1 0 62160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_551
timestamp 1663859327
transform 1 0 63056 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1663859327
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_562
timestamp 1663859327
transform 1 0 64288 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_594
timestamp 1663859327
transform 1 0 67872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1663859327
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_602
timestamp 1663859327
transform 1 0 68768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_608
timestamp 1663859327
transform 1 0 69440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_612
timestamp 1663859327
transform 1 0 69888 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_617
timestamp 1663859327
transform 1 0 70448 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_625
timestamp 1663859327
transform 1 0 71344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1663859327
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_632
timestamp 1663859327
transform 1 0 72128 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1663859327
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1663859327
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_672
timestamp 1663859327
transform 1 0 76608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_676
timestamp 1663859327
transform 1 0 77056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_678
timestamp 1663859327
transform 1 0 77280 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_683
timestamp 1663859327
transform 1 0 77840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_695
timestamp 1663859327
transform 1 0 79184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_699
timestamp 1663859327
transform 1 0 79632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_702
timestamp 1663859327
transform 1 0 79968 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_718
timestamp 1663859327
transform 1 0 81760 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_726
timestamp 1663859327
transform 1 0 82656 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_731
timestamp 1663859327
transform 1 0 83216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_737
timestamp 1663859327
transform 1 0 83888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_749
timestamp 1663859327
transform 1 0 85232 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_761
timestamp 1663859327
transform 1 0 86576 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_769
timestamp 1663859327
transform 1 0 87472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_772
timestamp 1663859327
transform 1 0 87808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_777
timestamp 1663859327
transform 1 0 88368 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_793
timestamp 1663859327
transform 1 0 90160 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_801
timestamp 1663859327
transform 1 0 91056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_807
timestamp 1663859327
transform 1 0 91728 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_827
timestamp 1663859327
transform 1 0 93968 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_835
timestamp 1663859327
transform 1 0 94864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_839
timestamp 1663859327
transform 1 0 95312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_842
timestamp 1663859327
transform 1 0 95648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1663859327
transform 1 0 99232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_877
timestamp 1663859327
transform 1 0 99568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_885
timestamp 1663859327
transform 1 0 100464 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_893
timestamp 1663859327
transform 1 0 101360 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_909
timestamp 1663859327
transform 1 0 103152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_912
timestamp 1663859327
transform 1 0 103488 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_944
timestamp 1663859327
transform 1 0 107072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_947
timestamp 1663859327
transform 1 0 107408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_952
timestamp 1663859327
transform 1 0 107968 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_960
timestamp 1663859327
transform 1 0 108864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_964
timestamp 1663859327
transform 1 0 109312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_966
timestamp 1663859327
transform 1 0 109536 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_971
timestamp 1663859327
transform 1 0 110096 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_979
timestamp 1663859327
transform 1 0 110992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1663859327
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_987
timestamp 1663859327
transform 1 0 111888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_995
timestamp 1663859327
transform 1 0 112784 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1011
timestamp 1663859327
transform 1 0 114576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1017
timestamp 1663859327
transform 1 0 115248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1025
timestamp 1663859327
transform 1 0 116144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1029
timestamp 1663859327
transform 1 0 116592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1044
timestamp 1663859327
transform 1 0 118272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1663859327
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_7 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2128 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1663859327
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1663859327
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1663859327
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1663859327
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1663859327
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1663859327
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1663859327
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1663859327
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1663859327
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1663859327
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1663859327
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1663859327
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1663859327
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1663859327
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1663859327
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_428
timestamp 1663859327
transform 1 0 49280 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1663859327
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1663859327
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_499
timestamp 1663859327
transform 1 0 57232 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_563
timestamp 1663859327
transform 1 0 64400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1663859327
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_570
timestamp 1663859327
transform 1 0 65184 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_634
timestamp 1663859327
transform 1 0 72352 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1663859327
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_641
timestamp 1663859327
transform 1 0 73136 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_705
timestamp 1663859327
transform 1 0 80304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_709
timestamp 1663859327
transform 1 0 80752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_712
timestamp 1663859327
transform 1 0 81088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_776
timestamp 1663859327
transform 1 0 88256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_780
timestamp 1663859327
transform 1 0 88704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_783
timestamp 1663859327
transform 1 0 89040 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_847
timestamp 1663859327
transform 1 0 96208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1663859327
transform 1 0 96656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_854
timestamp 1663859327
transform 1 0 96992 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_918
timestamp 1663859327
transform 1 0 104160 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_922
timestamp 1663859327
transform 1 0 104608 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_925
timestamp 1663859327
transform 1 0 104944 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_989
timestamp 1663859327
transform 1 0 112112 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_993
timestamp 1663859327
transform 1 0 112560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_996
timestamp 1663859327
transform 1 0 112896 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1030
timestamp 1663859327
transform 1 0 116704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1032
timestamp 1663859327
transform 1 0 116928 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1037
timestamp 1663859327
transform 1 0 117488 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1039
timestamp 1663859327
transform 1 0 117712 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1044
timestamp 1663859327
transform 1 0 118272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1663859327
transform 1 0 1568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_7
timestamp 1663859327
transform 1 0 2128 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_23
timestamp 1663859327
transform 1 0 3920 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_31
timestamp 1663859327
transform 1 0 4816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1663859327
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1663859327
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1663859327
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1663859327
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1663859327
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1663859327
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1663859327
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1663859327
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1663859327
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1663859327
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1663859327
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1663859327
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1663859327
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1663859327
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1663859327
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1663859327
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1663859327
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1663859327
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_463
timestamp 1663859327
transform 1 0 53200 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_527
timestamp 1663859327
transform 1 0 60368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1663859327
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_534
timestamp 1663859327
transform 1 0 61152 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_598
timestamp 1663859327
transform 1 0 68320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1663859327
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_605
timestamp 1663859327
transform 1 0 69104 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_669
timestamp 1663859327
transform 1 0 76272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1663859327
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_676
timestamp 1663859327
transform 1 0 77056 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_740
timestamp 1663859327
transform 1 0 84224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1663859327
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_747
timestamp 1663859327
transform 1 0 85008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_811
timestamp 1663859327
transform 1 0 92176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1663859327
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_818
timestamp 1663859327
transform 1 0 92960 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_882
timestamp 1663859327
transform 1 0 100128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_886
timestamp 1663859327
transform 1 0 100576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_889
timestamp 1663859327
transform 1 0 100912 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_953
timestamp 1663859327
transform 1 0 108080 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_957
timestamp 1663859327
transform 1 0 108528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_960
timestamp 1663859327
transform 1 0 108864 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1024
timestamp 1663859327
transform 1 0 116032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1028
timestamp 1663859327
transform 1 0 116480 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1031
timestamp 1663859327
transform 1 0 116816 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1039
timestamp 1663859327
transform 1 0 117712 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1044
timestamp 1663859327
transform 1 0 118272 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1663859327
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1663859327
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1663859327
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1663859327
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1663859327
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1663859327
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1663859327
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1663859327
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1663859327
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1663859327
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1663859327
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1663859327
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1663859327
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1663859327
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1663859327
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1663859327
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1663859327
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1663859327
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1663859327
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1663859327
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1663859327
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_499
timestamp 1663859327
transform 1 0 57232 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1663859327
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1663859327
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_570
timestamp 1663859327
transform 1 0 65184 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_634
timestamp 1663859327
transform 1 0 72352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1663859327
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_641
timestamp 1663859327
transform 1 0 73136 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_705
timestamp 1663859327
transform 1 0 80304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_709
timestamp 1663859327
transform 1 0 80752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_712
timestamp 1663859327
transform 1 0 81088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_776
timestamp 1663859327
transform 1 0 88256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_780
timestamp 1663859327
transform 1 0 88704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_783
timestamp 1663859327
transform 1 0 89040 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_847
timestamp 1663859327
transform 1 0 96208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_851
timestamp 1663859327
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_854
timestamp 1663859327
transform 1 0 96992 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_918
timestamp 1663859327
transform 1 0 104160 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_922
timestamp 1663859327
transform 1 0 104608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_925
timestamp 1663859327
transform 1 0 104944 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_989
timestamp 1663859327
transform 1 0 112112 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_993
timestamp 1663859327
transform 1 0 112560 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_996
timestamp 1663859327
transform 1 0 112896 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_1028
timestamp 1663859327
transform 1 0 116480 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1044
timestamp 1663859327
transform 1 0 118272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1663859327
transform 1 0 1568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_7
timestamp 1663859327
transform 1 0 2128 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_23
timestamp 1663859327
transform 1 0 3920 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_31
timestamp 1663859327
transform 1 0 4816 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1663859327
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1663859327
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1663859327
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1663859327
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1663859327
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1663859327
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1663859327
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1663859327
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1663859327
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1663859327
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1663859327
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1663859327
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1663859327
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1663859327
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1663859327
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1663859327
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1663859327
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1663859327
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1663859327
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1663859327
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1663859327
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1663859327
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_598
timestamp 1663859327
transform 1 0 68320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1663859327
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1663859327
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_669
timestamp 1663859327
transform 1 0 76272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1663859327
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_676
timestamp 1663859327
transform 1 0 77056 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_740
timestamp 1663859327
transform 1 0 84224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1663859327
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_747
timestamp 1663859327
transform 1 0 85008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_811
timestamp 1663859327
transform 1 0 92176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_815
timestamp 1663859327
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_818
timestamp 1663859327
transform 1 0 92960 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_882
timestamp 1663859327
transform 1 0 100128 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_886
timestamp 1663859327
transform 1 0 100576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_889
timestamp 1663859327
transform 1 0 100912 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_953
timestamp 1663859327
transform 1 0 108080 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_957
timestamp 1663859327
transform 1 0 108528 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_960
timestamp 1663859327
transform 1 0 108864 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1024
timestamp 1663859327
transform 1 0 116032 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1028
timestamp 1663859327
transform 1 0 116480 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1031
timestamp 1663859327
transform 1 0 116816 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1039
timestamp 1663859327
transform 1 0 117712 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1043
timestamp 1663859327
transform 1 0 118160 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1663859327
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1663859327
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1663859327
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1663859327
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1663859327
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1663859327
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1663859327
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1663859327
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1663859327
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1663859327
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1663859327
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1663859327
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1663859327
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1663859327
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1663859327
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1663859327
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1663859327
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1663859327
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1663859327
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1663859327
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1663859327
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1663859327
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1663859327
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1663859327
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1663859327
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1663859327
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1663859327
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_641
timestamp 1663859327
transform 1 0 73136 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_705
timestamp 1663859327
transform 1 0 80304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_709
timestamp 1663859327
transform 1 0 80752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_712
timestamp 1663859327
transform 1 0 81088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_776
timestamp 1663859327
transform 1 0 88256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1663859327
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_783
timestamp 1663859327
transform 1 0 89040 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_847
timestamp 1663859327
transform 1 0 96208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1663859327
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_854
timestamp 1663859327
transform 1 0 96992 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_918
timestamp 1663859327
transform 1 0 104160 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_922
timestamp 1663859327
transform 1 0 104608 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_925
timestamp 1663859327
transform 1 0 104944 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_989
timestamp 1663859327
transform 1 0 112112 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_993
timestamp 1663859327
transform 1 0 112560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_996
timestamp 1663859327
transform 1 0 112896 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_1028
timestamp 1663859327
transform 1 0 116480 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1044
timestamp 1663859327
transform 1 0 118272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1663859327
transform 1 0 1568 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_7
timestamp 1663859327
transform 1 0 2128 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_23
timestamp 1663859327
transform 1 0 3920 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_31
timestamp 1663859327
transform 1 0 4816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1663859327
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1663859327
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1663859327
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1663859327
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1663859327
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1663859327
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1663859327
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1663859327
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1663859327
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1663859327
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1663859327
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1663859327
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1663859327
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1663859327
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1663859327
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1663859327
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1663859327
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1663859327
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1663859327
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1663859327
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1663859327
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1663859327
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1663859327
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1663859327
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1663859327
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1663859327
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1663859327
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1663859327
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1663859327
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1663859327
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_747
timestamp 1663859327
transform 1 0 85008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_811
timestamp 1663859327
transform 1 0 92176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1663859327
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_818
timestamp 1663859327
transform 1 0 92960 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_882
timestamp 1663859327
transform 1 0 100128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1663859327
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_889
timestamp 1663859327
transform 1 0 100912 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_953
timestamp 1663859327
transform 1 0 108080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_957
timestamp 1663859327
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_960
timestamp 1663859327
transform 1 0 108864 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1024
timestamp 1663859327
transform 1 0 116032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1028
timestamp 1663859327
transform 1 0 116480 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1031
timestamp 1663859327
transform 1 0 116816 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1039
timestamp 1663859327
transform 1 0 117712 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1043
timestamp 1663859327
transform 1 0 118160 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1663859327
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1663859327
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1663859327
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1663859327
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1663859327
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1663859327
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1663859327
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1663859327
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1663859327
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1663859327
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1663859327
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1663859327
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1663859327
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1663859327
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1663859327
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1663859327
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1663859327
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1663859327
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1663859327
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1663859327
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1663859327
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1663859327
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1663859327
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1663859327
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1663859327
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1663859327
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1663859327
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1663859327
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1663859327
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1663859327
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1663859327
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1663859327
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1663859327
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_783
timestamp 1663859327
transform 1 0 89040 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_847
timestamp 1663859327
transform 1 0 96208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1663859327
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_854
timestamp 1663859327
transform 1 0 96992 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_918
timestamp 1663859327
transform 1 0 104160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1663859327
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_925
timestamp 1663859327
transform 1 0 104944 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_989
timestamp 1663859327
transform 1 0 112112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_993
timestamp 1663859327
transform 1 0 112560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_996
timestamp 1663859327
transform 1 0 112896 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_1028
timestamp 1663859327
transform 1 0 116480 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1044
timestamp 1663859327
transform 1 0 118272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1663859327
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1663859327
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1663859327
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1663859327
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1663859327
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1663859327
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1663859327
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1663859327
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1663859327
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1663859327
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1663859327
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1663859327
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1663859327
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1663859327
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1663859327
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1663859327
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1663859327
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1663859327
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1663859327
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1663859327
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1663859327
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1663859327
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1663859327
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1663859327
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1663859327
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1663859327
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1663859327
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1663859327
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1663859327
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1663859327
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1663859327
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1663859327
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1663859327
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1663859327
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1663859327
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_818
timestamp 1663859327
transform 1 0 92960 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_882
timestamp 1663859327
transform 1 0 100128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_886
timestamp 1663859327
transform 1 0 100576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_889
timestamp 1663859327
transform 1 0 100912 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_953
timestamp 1663859327
transform 1 0 108080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1663859327
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_960
timestamp 1663859327
transform 1 0 108864 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1024
timestamp 1663859327
transform 1 0 116032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1028
timestamp 1663859327
transform 1 0 116480 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_1031
timestamp 1663859327
transform 1 0 116816 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1039
timestamp 1663859327
transform 1 0 117712 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1043
timestamp 1663859327
transform 1 0 118160 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1663859327
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1663859327
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1663859327
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1663859327
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1663859327
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1663859327
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1663859327
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1663859327
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1663859327
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1663859327
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1663859327
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1663859327
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1663859327
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1663859327
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1663859327
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1663859327
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1663859327
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1663859327
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1663859327
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1663859327
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1663859327
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1663859327
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1663859327
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1663859327
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1663859327
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1663859327
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1663859327
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1663859327
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1663859327
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1663859327
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1663859327
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1663859327
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1663859327
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1663859327
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1663859327
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1663859327
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_854
timestamp 1663859327
transform 1 0 96992 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_918
timestamp 1663859327
transform 1 0 104160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1663859327
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_925
timestamp 1663859327
transform 1 0 104944 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_989
timestamp 1663859327
transform 1 0 112112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_993
timestamp 1663859327
transform 1 0 112560 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_996
timestamp 1663859327
transform 1 0 112896 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_1028
timestamp 1663859327
transform 1 0 116480 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1036
timestamp 1663859327
transform 1 0 117376 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1044
timestamp 1663859327
transform 1 0 118272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_2
timestamp 1663859327
transform 1 0 1568 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_7
timestamp 1663859327
transform 1 0 2128 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_23
timestamp 1663859327
transform 1 0 3920 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_31
timestamp 1663859327
transform 1 0 4816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1663859327
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1663859327
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1663859327
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1663859327
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1663859327
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1663859327
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1663859327
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1663859327
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1663859327
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1663859327
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1663859327
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1663859327
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1663859327
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1663859327
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1663859327
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1663859327
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1663859327
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1663859327
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1663859327
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1663859327
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1663859327
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1663859327
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1663859327
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1663859327
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1663859327
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1663859327
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1663859327
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1663859327
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1663859327
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1663859327
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1663859327
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1663859327
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1663859327
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_818
timestamp 1663859327
transform 1 0 92960 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_882
timestamp 1663859327
transform 1 0 100128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_886
timestamp 1663859327
transform 1 0 100576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_889
timestamp 1663859327
transform 1 0 100912 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_953
timestamp 1663859327
transform 1 0 108080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_957
timestamp 1663859327
transform 1 0 108528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_960
timestamp 1663859327
transform 1 0 108864 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1024
timestamp 1663859327
transform 1 0 116032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1663859327
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_1031
timestamp 1663859327
transform 1 0 116816 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1039
timestamp 1663859327
transform 1 0 117712 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1043
timestamp 1663859327
transform 1 0 118160 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1663859327
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1663859327
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1663859327
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1663859327
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1663859327
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1663859327
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1663859327
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1663859327
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1663859327
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1663859327
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1663859327
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1663859327
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1663859327
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1663859327
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1663859327
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1663859327
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1663859327
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1663859327
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1663859327
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1663859327
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1663859327
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1663859327
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1663859327
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1663859327
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1663859327
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1663859327
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1663859327
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1663859327
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1663859327
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1663859327
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1663859327
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1663859327
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1663859327
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1663859327
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1663859327
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1663859327
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_854
timestamp 1663859327
transform 1 0 96992 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_918
timestamp 1663859327
transform 1 0 104160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_922
timestamp 1663859327
transform 1 0 104608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_925
timestamp 1663859327
transform 1 0 104944 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_989
timestamp 1663859327
transform 1 0 112112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_993
timestamp 1663859327
transform 1 0 112560 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_996
timestamp 1663859327
transform 1 0 112896 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_1028
timestamp 1663859327
transform 1 0 116480 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1036
timestamp 1663859327
transform 1 0 117376 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1044
timestamp 1663859327
transform 1 0 118272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1663859327
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1663859327
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1663859327
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1663859327
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1663859327
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1663859327
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1663859327
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1663859327
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1663859327
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1663859327
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1663859327
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1663859327
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1663859327
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1663859327
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1663859327
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1663859327
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1663859327
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1663859327
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1663859327
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1663859327
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1663859327
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1663859327
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1663859327
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1663859327
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1663859327
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1663859327
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1663859327
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1663859327
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1663859327
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1663859327
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1663859327
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1663859327
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1663859327
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1663859327
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1663859327
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1663859327
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_882
timestamp 1663859327
transform 1 0 100128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1663859327
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_889
timestamp 1663859327
transform 1 0 100912 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_953
timestamp 1663859327
transform 1 0 108080 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_957
timestamp 1663859327
transform 1 0 108528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1663859327
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1663859327
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1663859327
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_1031
timestamp 1663859327
transform 1 0 116816 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1039
timestamp 1663859327
transform 1 0 117712 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_1043
timestamp 1663859327
transform 1 0 118160 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1663859327
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1663859327
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1663859327
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1663859327
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1663859327
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1663859327
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1663859327
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1663859327
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1663859327
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1663859327
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1663859327
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1663859327
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1663859327
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1663859327
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1663859327
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1663859327
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1663859327
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1663859327
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1663859327
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1663859327
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1663859327
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1663859327
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1663859327
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1663859327
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1663859327
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1663859327
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1663859327
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1663859327
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1663859327
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1663859327
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1663859327
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1663859327
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1663859327
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1663859327
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1663859327
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1663859327
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1663859327
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1663859327
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1663859327
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1663859327
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1663859327
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1663859327
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_996
timestamp 1663859327
transform 1 0 112896 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_1028
timestamp 1663859327
transform 1 0 116480 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1044
timestamp 1663859327
transform 1 0 118272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1663859327
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1663859327
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1663859327
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1663859327
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1663859327
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1663859327
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1663859327
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1663859327
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1663859327
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1663859327
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1663859327
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1663859327
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1663859327
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1663859327
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1663859327
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1663859327
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1663859327
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1663859327
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1663859327
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1663859327
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1663859327
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1663859327
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1663859327
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1663859327
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1663859327
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1663859327
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1663859327
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1663859327
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1663859327
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1663859327
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1663859327
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1663859327
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1663859327
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1663859327
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1663859327
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1663859327
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1663859327
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1663859327
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1663859327
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1663859327
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1663859327
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_960
timestamp 1663859327
transform 1 0 108864 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1024
timestamp 1663859327
transform 1 0 116032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1028
timestamp 1663859327
transform 1 0 116480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_1031
timestamp 1663859327
transform 1 0 116816 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1039
timestamp 1663859327
transform 1 0 117712 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1044
timestamp 1663859327
transform 1 0 118272 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1663859327
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1663859327
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1663859327
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1663859327
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1663859327
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1663859327
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1663859327
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1663859327
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1663859327
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1663859327
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1663859327
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1663859327
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1663859327
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1663859327
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1663859327
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1663859327
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1663859327
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1663859327
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1663859327
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1663859327
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1663859327
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1663859327
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1663859327
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1663859327
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1663859327
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1663859327
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1663859327
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1663859327
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1663859327
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1663859327
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1663859327
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1663859327
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1663859327
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1663859327
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1663859327
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1663859327
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1663859327
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1663859327
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1663859327
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1663859327
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1663859327
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1663859327
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_996
timestamp 1663859327
transform 1 0 112896 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_1028
timestamp 1663859327
transform 1 0 116480 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1044
timestamp 1663859327
transform 1 0 118272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1663859327
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1663859327
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1663859327
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1663859327
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1663859327
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1663859327
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1663859327
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1663859327
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1663859327
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1663859327
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1663859327
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1663859327
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1663859327
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1663859327
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1663859327
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1663859327
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1663859327
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1663859327
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1663859327
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1663859327
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1663859327
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1663859327
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1663859327
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1663859327
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1663859327
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1663859327
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1663859327
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1663859327
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1663859327
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_676
timestamp 1663859327
transform 1 0 77056 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_740
timestamp 1663859327
transform 1 0 84224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_744
timestamp 1663859327
transform 1 0 84672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_747
timestamp 1663859327
transform 1 0 85008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_811
timestamp 1663859327
transform 1 0 92176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_815
timestamp 1663859327
transform 1 0 92624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_818
timestamp 1663859327
transform 1 0 92960 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_882
timestamp 1663859327
transform 1 0 100128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_886
timestamp 1663859327
transform 1 0 100576 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_889
timestamp 1663859327
transform 1 0 100912 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_953
timestamp 1663859327
transform 1 0 108080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_957
timestamp 1663859327
transform 1 0 108528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_960
timestamp 1663859327
transform 1 0 108864 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1024
timestamp 1663859327
transform 1 0 116032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1028
timestamp 1663859327
transform 1 0 116480 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_1031
timestamp 1663859327
transform 1 0 116816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1039
timestamp 1663859327
transform 1 0 117712 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1043
timestamp 1663859327
transform 1 0 118160 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1663859327
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1663859327
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1663859327
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1663859327
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1663859327
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1663859327
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1663859327
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1663859327
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1663859327
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1663859327
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1663859327
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1663859327
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1663859327
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1663859327
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1663859327
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1663859327
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1663859327
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1663859327
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1663859327
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1663859327
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1663859327
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1663859327
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1663859327
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1663859327
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1663859327
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1663859327
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1663859327
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_641
timestamp 1663859327
transform 1 0 73136 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_705
timestamp 1663859327
transform 1 0 80304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_709
timestamp 1663859327
transform 1 0 80752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_712
timestamp 1663859327
transform 1 0 81088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_776
timestamp 1663859327
transform 1 0 88256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_780
timestamp 1663859327
transform 1 0 88704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_783
timestamp 1663859327
transform 1 0 89040 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_847
timestamp 1663859327
transform 1 0 96208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_851
timestamp 1663859327
transform 1 0 96656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_854
timestamp 1663859327
transform 1 0 96992 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_918
timestamp 1663859327
transform 1 0 104160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_922
timestamp 1663859327
transform 1 0 104608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_925
timestamp 1663859327
transform 1 0 104944 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_989
timestamp 1663859327
transform 1 0 112112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_993
timestamp 1663859327
transform 1 0 112560 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_996
timestamp 1663859327
transform 1 0 112896 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_1028
timestamp 1663859327
transform 1 0 116480 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1036
timestamp 1663859327
transform 1 0 117376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1044
timestamp 1663859327
transform 1 0 118272 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1663859327
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_7
timestamp 1663859327
transform 1 0 2128 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_23
timestamp 1663859327
transform 1 0 3920 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_31
timestamp 1663859327
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1663859327
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1663859327
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1663859327
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1663859327
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1663859327
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1663859327
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1663859327
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1663859327
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1663859327
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1663859327
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1663859327
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1663859327
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1663859327
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1663859327
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1663859327
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1663859327
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1663859327
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1663859327
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1663859327
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1663859327
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1663859327
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1663859327
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1663859327
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1663859327
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1663859327
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1663859327
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1663859327
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_676
timestamp 1663859327
transform 1 0 77056 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_740
timestamp 1663859327
transform 1 0 84224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_744
timestamp 1663859327
transform 1 0 84672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_747
timestamp 1663859327
transform 1 0 85008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_811
timestamp 1663859327
transform 1 0 92176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_815
timestamp 1663859327
transform 1 0 92624 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_818
timestamp 1663859327
transform 1 0 92960 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_882
timestamp 1663859327
transform 1 0 100128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_886
timestamp 1663859327
transform 1 0 100576 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_889
timestamp 1663859327
transform 1 0 100912 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_953
timestamp 1663859327
transform 1 0 108080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_957
timestamp 1663859327
transform 1 0 108528 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_960
timestamp 1663859327
transform 1 0 108864 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1024
timestamp 1663859327
transform 1 0 116032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1028
timestamp 1663859327
transform 1 0 116480 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_1031
timestamp 1663859327
transform 1 0 116816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1039
timestamp 1663859327
transform 1 0 117712 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1044
timestamp 1663859327
transform 1 0 118272 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1663859327
transform 1 0 1568 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_7
timestamp 1663859327
transform 1 0 2128 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1663859327
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1663859327
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1663859327
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1663859327
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1663859327
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1663859327
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1663859327
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1663859327
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1663859327
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1663859327
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1663859327
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1663859327
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1663859327
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1663859327
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1663859327
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1663859327
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1663859327
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1663859327
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1663859327
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1663859327
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1663859327
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1663859327
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1663859327
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1663859327
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_641
timestamp 1663859327
transform 1 0 73136 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_705
timestamp 1663859327
transform 1 0 80304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_709
timestamp 1663859327
transform 1 0 80752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_712
timestamp 1663859327
transform 1 0 81088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_776
timestamp 1663859327
transform 1 0 88256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_780
timestamp 1663859327
transform 1 0 88704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_783
timestamp 1663859327
transform 1 0 89040 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_847
timestamp 1663859327
transform 1 0 96208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_851
timestamp 1663859327
transform 1 0 96656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_854
timestamp 1663859327
transform 1 0 96992 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_918
timestamp 1663859327
transform 1 0 104160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_922
timestamp 1663859327
transform 1 0 104608 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_925
timestamp 1663859327
transform 1 0 104944 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_989
timestamp 1663859327
transform 1 0 112112 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_993
timestamp 1663859327
transform 1 0 112560 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_996
timestamp 1663859327
transform 1 0 112896 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_1028
timestamp 1663859327
transform 1 0 116480 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1044
timestamp 1663859327
transform 1 0 118272 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1663859327
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1663859327
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1663859327
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1663859327
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1663859327
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1663859327
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1663859327
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1663859327
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1663859327
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1663859327
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1663859327
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1663859327
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1663859327
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1663859327
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1663859327
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1663859327
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1663859327
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1663859327
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1663859327
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1663859327
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1663859327
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1663859327
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1663859327
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1663859327
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1663859327
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1663859327
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1663859327
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1663859327
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1663859327
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_676
timestamp 1663859327
transform 1 0 77056 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_740
timestamp 1663859327
transform 1 0 84224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_744
timestamp 1663859327
transform 1 0 84672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_747
timestamp 1663859327
transform 1 0 85008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_811
timestamp 1663859327
transform 1 0 92176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_815
timestamp 1663859327
transform 1 0 92624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_818
timestamp 1663859327
transform 1 0 92960 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_882
timestamp 1663859327
transform 1 0 100128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_886
timestamp 1663859327
transform 1 0 100576 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_889
timestamp 1663859327
transform 1 0 100912 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_953
timestamp 1663859327
transform 1 0 108080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_957
timestamp 1663859327
transform 1 0 108528 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_960
timestamp 1663859327
transform 1 0 108864 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1024
timestamp 1663859327
transform 1 0 116032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1028
timestamp 1663859327
transform 1 0 116480 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_1031
timestamp 1663859327
transform 1 0 116816 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1039
timestamp 1663859327
transform 1 0 117712 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_1043
timestamp 1663859327
transform 1 0 118160 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1663859327
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1663859327
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1663859327
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1663859327
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1663859327
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1663859327
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1663859327
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1663859327
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1663859327
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1663859327
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1663859327
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1663859327
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1663859327
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1663859327
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1663859327
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1663859327
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1663859327
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1663859327
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1663859327
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1663859327
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1663859327
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1663859327
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1663859327
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1663859327
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1663859327
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1663859327
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1663859327
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_641
timestamp 1663859327
transform 1 0 73136 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_705
timestamp 1663859327
transform 1 0 80304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_709
timestamp 1663859327
transform 1 0 80752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_712
timestamp 1663859327
transform 1 0 81088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_776
timestamp 1663859327
transform 1 0 88256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_780
timestamp 1663859327
transform 1 0 88704 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_783
timestamp 1663859327
transform 1 0 89040 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_847
timestamp 1663859327
transform 1 0 96208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_851
timestamp 1663859327
transform 1 0 96656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_854
timestamp 1663859327
transform 1 0 96992 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_918
timestamp 1663859327
transform 1 0 104160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_922
timestamp 1663859327
transform 1 0 104608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_925
timestamp 1663859327
transform 1 0 104944 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_989
timestamp 1663859327
transform 1 0 112112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_993
timestamp 1663859327
transform 1 0 112560 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_996
timestamp 1663859327
transform 1 0 112896 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_1028
timestamp 1663859327
transform 1 0 116480 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1044
timestamp 1663859327
transform 1 0 118272 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1663859327
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1663859327
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1663859327
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1663859327
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1663859327
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1663859327
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1663859327
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1663859327
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1663859327
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1663859327
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1663859327
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1663859327
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1663859327
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1663859327
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1663859327
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1663859327
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1663859327
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1663859327
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1663859327
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1663859327
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1663859327
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1663859327
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1663859327
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1663859327
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1663859327
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1663859327
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1663859327
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1663859327
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1663859327
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_676
timestamp 1663859327
transform 1 0 77056 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_740
timestamp 1663859327
transform 1 0 84224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_744
timestamp 1663859327
transform 1 0 84672 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_747
timestamp 1663859327
transform 1 0 85008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_811
timestamp 1663859327
transform 1 0 92176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_815
timestamp 1663859327
transform 1 0 92624 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_818
timestamp 1663859327
transform 1 0 92960 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_882
timestamp 1663859327
transform 1 0 100128 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_886
timestamp 1663859327
transform 1 0 100576 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_889
timestamp 1663859327
transform 1 0 100912 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_953
timestamp 1663859327
transform 1 0 108080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_957
timestamp 1663859327
transform 1 0 108528 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_960
timestamp 1663859327
transform 1 0 108864 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1024
timestamp 1663859327
transform 1 0 116032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1028
timestamp 1663859327
transform 1 0 116480 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_1031
timestamp 1663859327
transform 1 0 116816 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1039
timestamp 1663859327
transform 1 0 117712 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1044
timestamp 1663859327
transform 1 0 118272 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1663859327
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_7
timestamp 1663859327
transform 1 0 2128 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1663859327
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1663859327
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1663859327
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1663859327
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1663859327
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1663859327
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1663859327
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1663859327
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1663859327
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1663859327
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1663859327
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1663859327
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1663859327
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1663859327
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1663859327
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1663859327
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1663859327
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1663859327
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1663859327
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1663859327
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1663859327
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1663859327
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1663859327
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1663859327
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_641
timestamp 1663859327
transform 1 0 73136 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_705
timestamp 1663859327
transform 1 0 80304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_709
timestamp 1663859327
transform 1 0 80752 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_712
timestamp 1663859327
transform 1 0 81088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_776
timestamp 1663859327
transform 1 0 88256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_780
timestamp 1663859327
transform 1 0 88704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_783
timestamp 1663859327
transform 1 0 89040 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_847
timestamp 1663859327
transform 1 0 96208 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_851
timestamp 1663859327
transform 1 0 96656 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_854
timestamp 1663859327
transform 1 0 96992 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_918
timestamp 1663859327
transform 1 0 104160 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_922
timestamp 1663859327
transform 1 0 104608 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_925
timestamp 1663859327
transform 1 0 104944 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_989
timestamp 1663859327
transform 1 0 112112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_993
timestamp 1663859327
transform 1 0 112560 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_996
timestamp 1663859327
transform 1 0 112896 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_1028
timestamp 1663859327
transform 1 0 116480 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1044
timestamp 1663859327
transform 1 0 118272 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1663859327
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1663859327
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1663859327
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1663859327
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1663859327
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1663859327
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1663859327
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1663859327
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1663859327
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1663859327
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1663859327
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1663859327
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1663859327
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1663859327
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1663859327
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1663859327
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1663859327
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1663859327
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1663859327
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1663859327
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1663859327
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1663859327
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1663859327
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1663859327
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1663859327
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1663859327
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1663859327
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_669
timestamp 1663859327
transform 1 0 76272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1663859327
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_676
timestamp 1663859327
transform 1 0 77056 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_740
timestamp 1663859327
transform 1 0 84224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_744
timestamp 1663859327
transform 1 0 84672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_747
timestamp 1663859327
transform 1 0 85008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_811
timestamp 1663859327
transform 1 0 92176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_815
timestamp 1663859327
transform 1 0 92624 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_818
timestamp 1663859327
transform 1 0 92960 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_882
timestamp 1663859327
transform 1 0 100128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_886
timestamp 1663859327
transform 1 0 100576 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_889
timestamp 1663859327
transform 1 0 100912 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_953
timestamp 1663859327
transform 1 0 108080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_957
timestamp 1663859327
transform 1 0 108528 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_960
timestamp 1663859327
transform 1 0 108864 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1024
timestamp 1663859327
transform 1 0 116032 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1028
timestamp 1663859327
transform 1 0 116480 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_1031
timestamp 1663859327
transform 1 0 116816 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1039
timestamp 1663859327
transform 1 0 117712 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_1043
timestamp 1663859327
transform 1 0 118160 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1663859327
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_7
timestamp 1663859327
transform 1 0 2128 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1663859327
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1663859327
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1663859327
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1663859327
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1663859327
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1663859327
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1663859327
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1663859327
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1663859327
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1663859327
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1663859327
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1663859327
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1663859327
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1663859327
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1663859327
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1663859327
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1663859327
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1663859327
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1663859327
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1663859327
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1663859327
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1663859327
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1663859327
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1663859327
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_641
timestamp 1663859327
transform 1 0 73136 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_705
timestamp 1663859327
transform 1 0 80304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_709
timestamp 1663859327
transform 1 0 80752 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_712
timestamp 1663859327
transform 1 0 81088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_776
timestamp 1663859327
transform 1 0 88256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_780
timestamp 1663859327
transform 1 0 88704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_783
timestamp 1663859327
transform 1 0 89040 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_847
timestamp 1663859327
transform 1 0 96208 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_851
timestamp 1663859327
transform 1 0 96656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_854
timestamp 1663859327
transform 1 0 96992 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_918
timestamp 1663859327
transform 1 0 104160 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_922
timestamp 1663859327
transform 1 0 104608 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_925
timestamp 1663859327
transform 1 0 104944 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_989
timestamp 1663859327
transform 1 0 112112 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_993
timestamp 1663859327
transform 1 0 112560 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_996
timestamp 1663859327
transform 1 0 112896 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_1028
timestamp 1663859327
transform 1 0 116480 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1036
timestamp 1663859327
transform 1 0 117376 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1044
timestamp 1663859327
transform 1 0 118272 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1663859327
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1663859327
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1663859327
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1663859327
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1663859327
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1663859327
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1663859327
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1663859327
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1663859327
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1663859327
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1663859327
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1663859327
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1663859327
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1663859327
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1663859327
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1663859327
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1663859327
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1663859327
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1663859327
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1663859327
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1663859327
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1663859327
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1663859327
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1663859327
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1663859327
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1663859327
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1663859327
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1663859327
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1663859327
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_676
timestamp 1663859327
transform 1 0 77056 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_740
timestamp 1663859327
transform 1 0 84224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_744
timestamp 1663859327
transform 1 0 84672 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_747
timestamp 1663859327
transform 1 0 85008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_811
timestamp 1663859327
transform 1 0 92176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_815
timestamp 1663859327
transform 1 0 92624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_818
timestamp 1663859327
transform 1 0 92960 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_882
timestamp 1663859327
transform 1 0 100128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_886
timestamp 1663859327
transform 1 0 100576 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_889
timestamp 1663859327
transform 1 0 100912 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_953
timestamp 1663859327
transform 1 0 108080 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_957
timestamp 1663859327
transform 1 0 108528 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_960
timestamp 1663859327
transform 1 0 108864 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1024
timestamp 1663859327
transform 1 0 116032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1028
timestamp 1663859327
transform 1 0 116480 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_1031
timestamp 1663859327
transform 1 0 116816 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1039
timestamp 1663859327
transform 1 0 117712 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_1043
timestamp 1663859327
transform 1 0 118160 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1663859327
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1663859327
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1663859327
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1663859327
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1663859327
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1663859327
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1663859327
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1663859327
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1663859327
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1663859327
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1663859327
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1663859327
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1663859327
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1663859327
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1663859327
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1663859327
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1663859327
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1663859327
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1663859327
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1663859327
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1663859327
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1663859327
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1663859327
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1663859327
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1663859327
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1663859327
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1663859327
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_641
timestamp 1663859327
transform 1 0 73136 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_705
timestamp 1663859327
transform 1 0 80304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_709
timestamp 1663859327
transform 1 0 80752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_712
timestamp 1663859327
transform 1 0 81088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_776
timestamp 1663859327
transform 1 0 88256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_780
timestamp 1663859327
transform 1 0 88704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_783
timestamp 1663859327
transform 1 0 89040 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_847
timestamp 1663859327
transform 1 0 96208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_851
timestamp 1663859327
transform 1 0 96656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_854
timestamp 1663859327
transform 1 0 96992 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_918
timestamp 1663859327
transform 1 0 104160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_922
timestamp 1663859327
transform 1 0 104608 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_925
timestamp 1663859327
transform 1 0 104944 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_989
timestamp 1663859327
transform 1 0 112112 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_993
timestamp 1663859327
transform 1 0 112560 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_996
timestamp 1663859327
transform 1 0 112896 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_1028
timestamp 1663859327
transform 1 0 116480 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1044
timestamp 1663859327
transform 1 0 118272 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1663859327
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1663859327
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1663859327
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1663859327
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1663859327
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1663859327
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1663859327
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1663859327
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1663859327
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1663859327
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1663859327
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1663859327
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1663859327
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1663859327
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1663859327
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1663859327
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1663859327
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1663859327
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1663859327
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1663859327
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1663859327
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1663859327
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1663859327
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1663859327
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1663859327
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1663859327
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1663859327
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1663859327
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1663859327
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_676
timestamp 1663859327
transform 1 0 77056 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_740
timestamp 1663859327
transform 1 0 84224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_744
timestamp 1663859327
transform 1 0 84672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_747
timestamp 1663859327
transform 1 0 85008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_811
timestamp 1663859327
transform 1 0 92176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_815
timestamp 1663859327
transform 1 0 92624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_818
timestamp 1663859327
transform 1 0 92960 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_882
timestamp 1663859327
transform 1 0 100128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_886
timestamp 1663859327
transform 1 0 100576 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_889
timestamp 1663859327
transform 1 0 100912 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_953
timestamp 1663859327
transform 1 0 108080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_957
timestamp 1663859327
transform 1 0 108528 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_960
timestamp 1663859327
transform 1 0 108864 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1024
timestamp 1663859327
transform 1 0 116032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1028
timestamp 1663859327
transform 1 0 116480 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_1031
timestamp 1663859327
transform 1 0 116816 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1039
timestamp 1663859327
transform 1 0 117712 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1044
timestamp 1663859327
transform 1 0 118272 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_2
timestamp 1663859327
transform 1 0 1568 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_7
timestamp 1663859327
transform 1 0 2128 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1663859327
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1663859327
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1663859327
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1663859327
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1663859327
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1663859327
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1663859327
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1663859327
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1663859327
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1663859327
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1663859327
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1663859327
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1663859327
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1663859327
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1663859327
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1663859327
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1663859327
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1663859327
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1663859327
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1663859327
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1663859327
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1663859327
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1663859327
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1663859327
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_641
timestamp 1663859327
transform 1 0 73136 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_705
timestamp 1663859327
transform 1 0 80304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_709
timestamp 1663859327
transform 1 0 80752 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_712
timestamp 1663859327
transform 1 0 81088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_776
timestamp 1663859327
transform 1 0 88256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_780
timestamp 1663859327
transform 1 0 88704 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_783
timestamp 1663859327
transform 1 0 89040 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_847
timestamp 1663859327
transform 1 0 96208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_851
timestamp 1663859327
transform 1 0 96656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_854
timestamp 1663859327
transform 1 0 96992 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_918
timestamp 1663859327
transform 1 0 104160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_922
timestamp 1663859327
transform 1 0 104608 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_925
timestamp 1663859327
transform 1 0 104944 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_989
timestamp 1663859327
transform 1 0 112112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_993
timestamp 1663859327
transform 1 0 112560 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_996
timestamp 1663859327
transform 1 0 112896 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_1028
timestamp 1663859327
transform 1 0 116480 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1044
timestamp 1663859327
transform 1 0 118272 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1663859327
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1663859327
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1663859327
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1663859327
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1663859327
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1663859327
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1663859327
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1663859327
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1663859327
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1663859327
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1663859327
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1663859327
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1663859327
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1663859327
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1663859327
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1663859327
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1663859327
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1663859327
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1663859327
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1663859327
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1663859327
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1663859327
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1663859327
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1663859327
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1663859327
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1663859327
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1663859327
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1663859327
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1663859327
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_676
timestamp 1663859327
transform 1 0 77056 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_740
timestamp 1663859327
transform 1 0 84224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_744
timestamp 1663859327
transform 1 0 84672 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_747
timestamp 1663859327
transform 1 0 85008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_811
timestamp 1663859327
transform 1 0 92176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_815
timestamp 1663859327
transform 1 0 92624 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_818
timestamp 1663859327
transform 1 0 92960 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_882
timestamp 1663859327
transform 1 0 100128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_886
timestamp 1663859327
transform 1 0 100576 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_889
timestamp 1663859327
transform 1 0 100912 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_953
timestamp 1663859327
transform 1 0 108080 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_957
timestamp 1663859327
transform 1 0 108528 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_960
timestamp 1663859327
transform 1 0 108864 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1024
timestamp 1663859327
transform 1 0 116032 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1028
timestamp 1663859327
transform 1 0 116480 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_1031
timestamp 1663859327
transform 1 0 116816 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1039
timestamp 1663859327
transform 1 0 117712 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1044
timestamp 1663859327
transform 1 0 118272 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1663859327
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1663859327
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1663859327
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1663859327
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1663859327
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1663859327
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1663859327
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1663859327
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1663859327
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1663859327
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1663859327
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1663859327
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1663859327
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1663859327
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1663859327
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1663859327
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1663859327
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1663859327
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1663859327
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1663859327
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1663859327
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1663859327
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1663859327
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1663859327
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1663859327
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1663859327
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1663859327
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_641
timestamp 1663859327
transform 1 0 73136 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_705
timestamp 1663859327
transform 1 0 80304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_709
timestamp 1663859327
transform 1 0 80752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_712
timestamp 1663859327
transform 1 0 81088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_776
timestamp 1663859327
transform 1 0 88256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_780
timestamp 1663859327
transform 1 0 88704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_783
timestamp 1663859327
transform 1 0 89040 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_847
timestamp 1663859327
transform 1 0 96208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_851
timestamp 1663859327
transform 1 0 96656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_854
timestamp 1663859327
transform 1 0 96992 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_918
timestamp 1663859327
transform 1 0 104160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_922
timestamp 1663859327
transform 1 0 104608 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_925
timestamp 1663859327
transform 1 0 104944 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_989
timestamp 1663859327
transform 1 0 112112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_993
timestamp 1663859327
transform 1 0 112560 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_996
timestamp 1663859327
transform 1 0 112896 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_1028
timestamp 1663859327
transform 1 0 116480 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1044
timestamp 1663859327
transform 1 0 118272 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1663859327
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1663859327
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1663859327
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1663859327
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1663859327
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1663859327
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1663859327
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1663859327
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1663859327
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1663859327
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1663859327
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1663859327
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1663859327
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1663859327
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1663859327
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1663859327
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1663859327
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1663859327
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1663859327
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1663859327
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1663859327
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1663859327
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1663859327
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1663859327
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1663859327
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1663859327
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1663859327
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1663859327
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1663859327
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_676
timestamp 1663859327
transform 1 0 77056 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_740
timestamp 1663859327
transform 1 0 84224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_744
timestamp 1663859327
transform 1 0 84672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_747
timestamp 1663859327
transform 1 0 85008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_811
timestamp 1663859327
transform 1 0 92176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_815
timestamp 1663859327
transform 1 0 92624 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_818
timestamp 1663859327
transform 1 0 92960 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_882
timestamp 1663859327
transform 1 0 100128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_886
timestamp 1663859327
transform 1 0 100576 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_889
timestamp 1663859327
transform 1 0 100912 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_953
timestamp 1663859327
transform 1 0 108080 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_957
timestamp 1663859327
transform 1 0 108528 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_960
timestamp 1663859327
transform 1 0 108864 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1024
timestamp 1663859327
transform 1 0 116032 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1028
timestamp 1663859327
transform 1 0 116480 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_1031
timestamp 1663859327
transform 1 0 116816 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1039
timestamp 1663859327
transform 1 0 117712 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_1043
timestamp 1663859327
transform 1 0 118160 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1663859327
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1663859327
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1663859327
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1663859327
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1663859327
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1663859327
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1663859327
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1663859327
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1663859327
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1663859327
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1663859327
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1663859327
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1663859327
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1663859327
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1663859327
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1663859327
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1663859327
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1663859327
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1663859327
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1663859327
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1663859327
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1663859327
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1663859327
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1663859327
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1663859327
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1663859327
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1663859327
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_641
timestamp 1663859327
transform 1 0 73136 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_705
timestamp 1663859327
transform 1 0 80304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_709
timestamp 1663859327
transform 1 0 80752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_712
timestamp 1663859327
transform 1 0 81088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_776
timestamp 1663859327
transform 1 0 88256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_780
timestamp 1663859327
transform 1 0 88704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_783
timestamp 1663859327
transform 1 0 89040 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_847
timestamp 1663859327
transform 1 0 96208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_851
timestamp 1663859327
transform 1 0 96656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_854
timestamp 1663859327
transform 1 0 96992 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_918
timestamp 1663859327
transform 1 0 104160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_922
timestamp 1663859327
transform 1 0 104608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_925
timestamp 1663859327
transform 1 0 104944 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_989
timestamp 1663859327
transform 1 0 112112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_993
timestamp 1663859327
transform 1 0 112560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_996
timestamp 1663859327
transform 1 0 112896 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_1028
timestamp 1663859327
transform 1 0 116480 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1036
timestamp 1663859327
transform 1 0 117376 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1044
timestamp 1663859327
transform 1 0 118272 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1663859327
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_7
timestamp 1663859327
transform 1 0 2128 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_23
timestamp 1663859327
transform 1 0 3920 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_31
timestamp 1663859327
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1663859327
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1663859327
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1663859327
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1663859327
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1663859327
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1663859327
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1663859327
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1663859327
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1663859327
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1663859327
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1663859327
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1663859327
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1663859327
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1663859327
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1663859327
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1663859327
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1663859327
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1663859327
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1663859327
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1663859327
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1663859327
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1663859327
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1663859327
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1663859327
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1663859327
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1663859327
transform 1 0 76272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1663859327
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_676
timestamp 1663859327
transform 1 0 77056 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_740
timestamp 1663859327
transform 1 0 84224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_744
timestamp 1663859327
transform 1 0 84672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_747
timestamp 1663859327
transform 1 0 85008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_811
timestamp 1663859327
transform 1 0 92176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_815
timestamp 1663859327
transform 1 0 92624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_818
timestamp 1663859327
transform 1 0 92960 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_882
timestamp 1663859327
transform 1 0 100128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_886
timestamp 1663859327
transform 1 0 100576 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_889
timestamp 1663859327
transform 1 0 100912 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_953
timestamp 1663859327
transform 1 0 108080 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_957
timestamp 1663859327
transform 1 0 108528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_960
timestamp 1663859327
transform 1 0 108864 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1024
timestamp 1663859327
transform 1 0 116032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1028
timestamp 1663859327
transform 1 0 116480 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_1031
timestamp 1663859327
transform 1 0 116816 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1039
timestamp 1663859327
transform 1 0 117712 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_1043
timestamp 1663859327
transform 1 0 118160 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1663859327
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1663859327
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1663859327
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1663859327
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1663859327
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1663859327
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1663859327
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1663859327
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1663859327
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1663859327
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1663859327
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1663859327
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1663859327
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1663859327
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1663859327
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1663859327
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1663859327
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1663859327
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1663859327
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1663859327
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1663859327
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1663859327
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1663859327
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1663859327
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1663859327
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1663859327
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1663859327
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_641
timestamp 1663859327
transform 1 0 73136 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_705
timestamp 1663859327
transform 1 0 80304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_709
timestamp 1663859327
transform 1 0 80752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_712
timestamp 1663859327
transform 1 0 81088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_776
timestamp 1663859327
transform 1 0 88256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_780
timestamp 1663859327
transform 1 0 88704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_783
timestamp 1663859327
transform 1 0 89040 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_847
timestamp 1663859327
transform 1 0 96208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_851
timestamp 1663859327
transform 1 0 96656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_854
timestamp 1663859327
transform 1 0 96992 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_918
timestamp 1663859327
transform 1 0 104160 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_922
timestamp 1663859327
transform 1 0 104608 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_925
timestamp 1663859327
transform 1 0 104944 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_989
timestamp 1663859327
transform 1 0 112112 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_993
timestamp 1663859327
transform 1 0 112560 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_996
timestamp 1663859327
transform 1 0 112896 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_1028
timestamp 1663859327
transform 1 0 116480 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1044
timestamp 1663859327
transform 1 0 118272 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1663859327
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1663859327
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1663859327
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1663859327
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1663859327
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1663859327
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1663859327
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1663859327
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1663859327
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1663859327
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1663859327
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1663859327
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1663859327
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1663859327
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1663859327
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1663859327
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1663859327
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1663859327
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1663859327
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1663859327
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1663859327
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1663859327
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1663859327
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1663859327
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1663859327
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1663859327
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1663859327
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1663859327
transform 1 0 76272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1663859327
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_676
timestamp 1663859327
transform 1 0 77056 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_740
timestamp 1663859327
transform 1 0 84224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_744
timestamp 1663859327
transform 1 0 84672 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_747
timestamp 1663859327
transform 1 0 85008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_811
timestamp 1663859327
transform 1 0 92176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_815
timestamp 1663859327
transform 1 0 92624 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_818
timestamp 1663859327
transform 1 0 92960 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_882
timestamp 1663859327
transform 1 0 100128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_886
timestamp 1663859327
transform 1 0 100576 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_889
timestamp 1663859327
transform 1 0 100912 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_953
timestamp 1663859327
transform 1 0 108080 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_957
timestamp 1663859327
transform 1 0 108528 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_960
timestamp 1663859327
transform 1 0 108864 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1024
timestamp 1663859327
transform 1 0 116032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1028
timestamp 1663859327
transform 1 0 116480 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_1031
timestamp 1663859327
transform 1 0 116816 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1039
timestamp 1663859327
transform 1 0 117712 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1044
timestamp 1663859327
transform 1 0 118272 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1663859327
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1663859327
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1663859327
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1663859327
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1663859327
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1663859327
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1663859327
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1663859327
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1663859327
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1663859327
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1663859327
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1663859327
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1663859327
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1663859327
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1663859327
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1663859327
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1663859327
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1663859327
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1663859327
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1663859327
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1663859327
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1663859327
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1663859327
transform 1 0 64400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1663859327
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1663859327
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1663859327
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1663859327
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_641
timestamp 1663859327
transform 1 0 73136 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_705
timestamp 1663859327
transform 1 0 80304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_709
timestamp 1663859327
transform 1 0 80752 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_712
timestamp 1663859327
transform 1 0 81088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_776
timestamp 1663859327
transform 1 0 88256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_780
timestamp 1663859327
transform 1 0 88704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_783
timestamp 1663859327
transform 1 0 89040 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_847
timestamp 1663859327
transform 1 0 96208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_851
timestamp 1663859327
transform 1 0 96656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_854
timestamp 1663859327
transform 1 0 96992 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_918
timestamp 1663859327
transform 1 0 104160 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_922
timestamp 1663859327
transform 1 0 104608 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_925
timestamp 1663859327
transform 1 0 104944 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_989
timestamp 1663859327
transform 1 0 112112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_993
timestamp 1663859327
transform 1 0 112560 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_996
timestamp 1663859327
transform 1 0 112896 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_1028
timestamp 1663859327
transform 1 0 116480 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1044
timestamp 1663859327
transform 1 0 118272 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1663859327
transform 1 0 1568 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_7
timestamp 1663859327
transform 1 0 2128 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_23
timestamp 1663859327
transform 1 0 3920 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_31
timestamp 1663859327
transform 1 0 4816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1663859327
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1663859327
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1663859327
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1663859327
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1663859327
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1663859327
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1663859327
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1663859327
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1663859327
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1663859327
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1663859327
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1663859327
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1663859327
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1663859327
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1663859327
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1663859327
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1663859327
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1663859327
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1663859327
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1663859327
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1663859327
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1663859327
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1663859327
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1663859327
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1663859327
transform 1 0 69104 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_669
timestamp 1663859327
transform 1 0 76272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1663859327
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_676
timestamp 1663859327
transform 1 0 77056 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_740
timestamp 1663859327
transform 1 0 84224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_744
timestamp 1663859327
transform 1 0 84672 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_747
timestamp 1663859327
transform 1 0 85008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_811
timestamp 1663859327
transform 1 0 92176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_815
timestamp 1663859327
transform 1 0 92624 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_818
timestamp 1663859327
transform 1 0 92960 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_882
timestamp 1663859327
transform 1 0 100128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_886
timestamp 1663859327
transform 1 0 100576 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_889
timestamp 1663859327
transform 1 0 100912 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_953
timestamp 1663859327
transform 1 0 108080 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_957
timestamp 1663859327
transform 1 0 108528 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_960
timestamp 1663859327
transform 1 0 108864 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1024
timestamp 1663859327
transform 1 0 116032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1028
timestamp 1663859327
transform 1 0 116480 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_1031
timestamp 1663859327
transform 1 0 116816 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1039
timestamp 1663859327
transform 1 0 117712 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1043
timestamp 1663859327
transform 1 0 118160 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1663859327
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1663859327
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1663859327
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1663859327
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1663859327
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1663859327
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1663859327
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1663859327
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1663859327
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1663859327
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1663859327
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1663859327
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1663859327
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1663859327
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1663859327
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1663859327
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1663859327
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1663859327
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1663859327
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1663859327
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1663859327
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1663859327
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1663859327
transform 1 0 64400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1663859327
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1663859327
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1663859327
transform 1 0 72352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1663859327
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_641
timestamp 1663859327
transform 1 0 73136 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_705
timestamp 1663859327
transform 1 0 80304 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_709
timestamp 1663859327
transform 1 0 80752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_712
timestamp 1663859327
transform 1 0 81088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_776
timestamp 1663859327
transform 1 0 88256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_780
timestamp 1663859327
transform 1 0 88704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_783
timestamp 1663859327
transform 1 0 89040 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_847
timestamp 1663859327
transform 1 0 96208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_851
timestamp 1663859327
transform 1 0 96656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_854
timestamp 1663859327
transform 1 0 96992 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_918
timestamp 1663859327
transform 1 0 104160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_922
timestamp 1663859327
transform 1 0 104608 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_925
timestamp 1663859327
transform 1 0 104944 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_989
timestamp 1663859327
transform 1 0 112112 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_993
timestamp 1663859327
transform 1 0 112560 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_996
timestamp 1663859327
transform 1 0 112896 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_1028
timestamp 1663859327
transform 1 0 116480 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1044
timestamp 1663859327
transform 1 0 118272 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1663859327
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1663859327
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1663859327
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1663859327
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1663859327
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1663859327
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1663859327
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1663859327
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1663859327
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1663859327
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1663859327
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1663859327
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1663859327
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1663859327
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1663859327
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1663859327
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1663859327
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1663859327
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1663859327
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1663859327
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1663859327
transform 1 0 53200 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1663859327
transform 1 0 60368 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1663859327
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1663859327
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1663859327
transform 1 0 68320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1663859327
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1663859327
transform 1 0 69104 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_669
timestamp 1663859327
transform 1 0 76272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1663859327
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_676
timestamp 1663859327
transform 1 0 77056 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_740
timestamp 1663859327
transform 1 0 84224 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_744
timestamp 1663859327
transform 1 0 84672 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_747
timestamp 1663859327
transform 1 0 85008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_811
timestamp 1663859327
transform 1 0 92176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_815
timestamp 1663859327
transform 1 0 92624 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_818
timestamp 1663859327
transform 1 0 92960 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_882
timestamp 1663859327
transform 1 0 100128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_886
timestamp 1663859327
transform 1 0 100576 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_889
timestamp 1663859327
transform 1 0 100912 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_953
timestamp 1663859327
transform 1 0 108080 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_957
timestamp 1663859327
transform 1 0 108528 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_960
timestamp 1663859327
transform 1 0 108864 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1024
timestamp 1663859327
transform 1 0 116032 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1028
timestamp 1663859327
transform 1 0 116480 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_1031
timestamp 1663859327
transform 1 0 116816 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1039
timestamp 1663859327
transform 1 0 117712 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1043
timestamp 1663859327
transform 1 0 118160 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1663859327
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1663859327
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1663859327
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1663859327
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1663859327
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1663859327
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1663859327
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1663859327
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1663859327
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1663859327
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1663859327
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1663859327
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1663859327
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1663859327
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1663859327
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1663859327
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1663859327
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1663859327
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1663859327
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1663859327
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1663859327
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1663859327
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1663859327
transform 1 0 64400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1663859327
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1663859327
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1663859327
transform 1 0 72352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1663859327
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_641
timestamp 1663859327
transform 1 0 73136 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_705
timestamp 1663859327
transform 1 0 80304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_709
timestamp 1663859327
transform 1 0 80752 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_712
timestamp 1663859327
transform 1 0 81088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_776
timestamp 1663859327
transform 1 0 88256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_780
timestamp 1663859327
transform 1 0 88704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_783
timestamp 1663859327
transform 1 0 89040 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_847
timestamp 1663859327
transform 1 0 96208 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_851
timestamp 1663859327
transform 1 0 96656 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_854
timestamp 1663859327
transform 1 0 96992 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_918
timestamp 1663859327
transform 1 0 104160 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_922
timestamp 1663859327
transform 1 0 104608 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_925
timestamp 1663859327
transform 1 0 104944 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_989
timestamp 1663859327
transform 1 0 112112 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_993
timestamp 1663859327
transform 1 0 112560 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_996
timestamp 1663859327
transform 1 0 112896 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_1012
timestamp 1663859327
transform 1 0 114688 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1020
timestamp 1663859327
transform 1 0 115584 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1024
timestamp 1663859327
transform 1 0 116032 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1028
timestamp 1663859327
transform 1 0 116480 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1044
timestamp 1663859327
transform 1 0 118272 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1663859327
transform 1 0 1568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_7
timestamp 1663859327
transform 1 0 2128 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_23
timestamp 1663859327
transform 1 0 3920 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_31
timestamp 1663859327
transform 1 0 4816 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1663859327
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1663859327
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1663859327
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1663859327
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1663859327
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1663859327
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1663859327
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1663859327
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1663859327
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1663859327
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1663859327
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1663859327
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1663859327
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1663859327
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1663859327
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1663859327
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_456
timestamp 1663859327
transform 1 0 52416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1663859327
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_463
timestamp 1663859327
transform 1 0 53200 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_527
timestamp 1663859327
transform 1 0 60368 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_531
timestamp 1663859327
transform 1 0 60816 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_534
timestamp 1663859327
transform 1 0 61152 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_598
timestamp 1663859327
transform 1 0 68320 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_602
timestamp 1663859327
transform 1 0 68768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_605
timestamp 1663859327
transform 1 0 69104 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_669
timestamp 1663859327
transform 1 0 76272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_673
timestamp 1663859327
transform 1 0 76720 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_676
timestamp 1663859327
transform 1 0 77056 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_740
timestamp 1663859327
transform 1 0 84224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_744
timestamp 1663859327
transform 1 0 84672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_747
timestamp 1663859327
transform 1 0 85008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_811
timestamp 1663859327
transform 1 0 92176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_815
timestamp 1663859327
transform 1 0 92624 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_818
timestamp 1663859327
transform 1 0 92960 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_882
timestamp 1663859327
transform 1 0 100128 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_886
timestamp 1663859327
transform 1 0 100576 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_889
timestamp 1663859327
transform 1 0 100912 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_953
timestamp 1663859327
transform 1 0 108080 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_957
timestamp 1663859327
transform 1 0 108528 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_960
timestamp 1663859327
transform 1 0 108864 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1024
timestamp 1663859327
transform 1 0 116032 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1028
timestamp 1663859327
transform 1 0 116480 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_1031
timestamp 1663859327
transform 1 0 116816 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1039
timestamp 1663859327
transform 1 0 117712 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1043
timestamp 1663859327
transform 1 0 118160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1663859327
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_7
timestamp 1663859327
transform 1 0 2128 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1663859327
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1663859327
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1663859327
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1663859327
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1663859327
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1663859327
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1663859327
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1663859327
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1663859327
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1663859327
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1663859327
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1663859327
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1663859327
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1663859327
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1663859327
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_428
timestamp 1663859327
transform 1 0 49280 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_492
timestamp 1663859327
transform 1 0 56448 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1663859327
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_499
timestamp 1663859327
transform 1 0 57232 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_563
timestamp 1663859327
transform 1 0 64400 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_567
timestamp 1663859327
transform 1 0 64848 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_570
timestamp 1663859327
transform 1 0 65184 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_634
timestamp 1663859327
transform 1 0 72352 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_638
timestamp 1663859327
transform 1 0 72800 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_641
timestamp 1663859327
transform 1 0 73136 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_705
timestamp 1663859327
transform 1 0 80304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_709
timestamp 1663859327
transform 1 0 80752 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_712
timestamp 1663859327
transform 1 0 81088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_776
timestamp 1663859327
transform 1 0 88256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_780
timestamp 1663859327
transform 1 0 88704 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_783
timestamp 1663859327
transform 1 0 89040 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_847
timestamp 1663859327
transform 1 0 96208 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_851
timestamp 1663859327
transform 1 0 96656 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_854
timestamp 1663859327
transform 1 0 96992 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_918
timestamp 1663859327
transform 1 0 104160 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_922
timestamp 1663859327
transform 1 0 104608 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_925
timestamp 1663859327
transform 1 0 104944 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_989
timestamp 1663859327
transform 1 0 112112 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_993
timestamp 1663859327
transform 1 0 112560 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_996
timestamp 1663859327
transform 1 0 112896 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_1028
timestamp 1663859327
transform 1 0 116480 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_1044
timestamp 1663859327
transform 1 0 118272 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1663859327
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1663859327
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1663859327
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1663859327
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1663859327
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1663859327
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1663859327
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1663859327
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1663859327
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1663859327
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1663859327
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1663859327
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1663859327
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1663859327
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1663859327
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1663859327
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1663859327
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1663859327
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1663859327
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1663859327
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_463
timestamp 1663859327
transform 1 0 53200 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_527
timestamp 1663859327
transform 1 0 60368 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_531
timestamp 1663859327
transform 1 0 60816 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_534
timestamp 1663859327
transform 1 0 61152 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_598
timestamp 1663859327
transform 1 0 68320 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_602
timestamp 1663859327
transform 1 0 68768 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_605
timestamp 1663859327
transform 1 0 69104 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_669
timestamp 1663859327
transform 1 0 76272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_673
timestamp 1663859327
transform 1 0 76720 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_676
timestamp 1663859327
transform 1 0 77056 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_740
timestamp 1663859327
transform 1 0 84224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_744
timestamp 1663859327
transform 1 0 84672 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_747
timestamp 1663859327
transform 1 0 85008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_811
timestamp 1663859327
transform 1 0 92176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_815
timestamp 1663859327
transform 1 0 92624 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_818
timestamp 1663859327
transform 1 0 92960 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_882
timestamp 1663859327
transform 1 0 100128 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_886
timestamp 1663859327
transform 1 0 100576 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_889
timestamp 1663859327
transform 1 0 100912 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_953
timestamp 1663859327
transform 1 0 108080 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_957
timestamp 1663859327
transform 1 0 108528 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_960
timestamp 1663859327
transform 1 0 108864 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1024
timestamp 1663859327
transform 1 0 116032 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_1028
timestamp 1663859327
transform 1 0 116480 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_1031
timestamp 1663859327
transform 1 0 116816 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_1039
timestamp 1663859327
transform 1 0 117712 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_1043
timestamp 1663859327
transform 1 0 118160 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1663859327
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1663859327
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1663859327
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1663859327
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1663859327
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1663859327
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1663859327
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1663859327
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1663859327
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1663859327
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1663859327
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1663859327
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1663859327
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1663859327
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1663859327
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1663859327
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1663859327
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1663859327
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_428
timestamp 1663859327
transform 1 0 49280 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_492
timestamp 1663859327
transform 1 0 56448 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1663859327
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_499
timestamp 1663859327
transform 1 0 57232 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_563
timestamp 1663859327
transform 1 0 64400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_567
timestamp 1663859327
transform 1 0 64848 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_570
timestamp 1663859327
transform 1 0 65184 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_634
timestamp 1663859327
transform 1 0 72352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_638
timestamp 1663859327
transform 1 0 72800 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_641
timestamp 1663859327
transform 1 0 73136 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_705
timestamp 1663859327
transform 1 0 80304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_709
timestamp 1663859327
transform 1 0 80752 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_712
timestamp 1663859327
transform 1 0 81088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_776
timestamp 1663859327
transform 1 0 88256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_780
timestamp 1663859327
transform 1 0 88704 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_783
timestamp 1663859327
transform 1 0 89040 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_847
timestamp 1663859327
transform 1 0 96208 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_851
timestamp 1663859327
transform 1 0 96656 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_854
timestamp 1663859327
transform 1 0 96992 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_918
timestamp 1663859327
transform 1 0 104160 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_922
timestamp 1663859327
transform 1 0 104608 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_925
timestamp 1663859327
transform 1 0 104944 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_989
timestamp 1663859327
transform 1 0 112112 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_993
timestamp 1663859327
transform 1 0 112560 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_996
timestamp 1663859327
transform 1 0 112896 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_1028
timestamp 1663859327
transform 1 0 116480 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_1036
timestamp 1663859327
transform 1 0 117376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_1044
timestamp 1663859327
transform 1 0 118272 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_2
timestamp 1663859327
transform 1 0 1568 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_7
timestamp 1663859327
transform 1 0 2128 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_23
timestamp 1663859327
transform 1 0 3920 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_31
timestamp 1663859327
transform 1 0 4816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1663859327
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1663859327
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1663859327
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1663859327
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1663859327
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1663859327
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1663859327
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1663859327
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1663859327
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1663859327
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1663859327
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1663859327
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1663859327
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1663859327
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1663859327
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_392
timestamp 1663859327
transform 1 0 45248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_456
timestamp 1663859327
transform 1 0 52416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1663859327
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_463
timestamp 1663859327
transform 1 0 53200 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_527
timestamp 1663859327
transform 1 0 60368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_531
timestamp 1663859327
transform 1 0 60816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_534
timestamp 1663859327
transform 1 0 61152 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_598
timestamp 1663859327
transform 1 0 68320 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_602
timestamp 1663859327
transform 1 0 68768 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_605
timestamp 1663859327
transform 1 0 69104 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_669
timestamp 1663859327
transform 1 0 76272 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_673
timestamp 1663859327
transform 1 0 76720 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_676
timestamp 1663859327
transform 1 0 77056 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_740
timestamp 1663859327
transform 1 0 84224 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_744
timestamp 1663859327
transform 1 0 84672 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_747
timestamp 1663859327
transform 1 0 85008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_811
timestamp 1663859327
transform 1 0 92176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_815
timestamp 1663859327
transform 1 0 92624 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_818
timestamp 1663859327
transform 1 0 92960 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_882
timestamp 1663859327
transform 1 0 100128 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_886
timestamp 1663859327
transform 1 0 100576 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_889
timestamp 1663859327
transform 1 0 100912 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_953
timestamp 1663859327
transform 1 0 108080 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_957
timestamp 1663859327
transform 1 0 108528 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_960
timestamp 1663859327
transform 1 0 108864 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1024
timestamp 1663859327
transform 1 0 116032 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_1028
timestamp 1663859327
transform 1 0 116480 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_1031
timestamp 1663859327
transform 1 0 116816 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_1039
timestamp 1663859327
transform 1 0 117712 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_1043
timestamp 1663859327
transform 1 0 118160 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1663859327
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1663859327
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1663859327
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1663859327
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1663859327
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1663859327
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1663859327
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1663859327
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1663859327
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1663859327
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1663859327
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1663859327
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1663859327
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1663859327
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1663859327
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_357
timestamp 1663859327
transform 1 0 41328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_421
timestamp 1663859327
transform 1 0 48496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_425
timestamp 1663859327
transform 1 0 48944 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1663859327
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1663859327
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1663859327
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_499
timestamp 1663859327
transform 1 0 57232 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_563
timestamp 1663859327
transform 1 0 64400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_567
timestamp 1663859327
transform 1 0 64848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_570
timestamp 1663859327
transform 1 0 65184 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_634
timestamp 1663859327
transform 1 0 72352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_638
timestamp 1663859327
transform 1 0 72800 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_641
timestamp 1663859327
transform 1 0 73136 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_705
timestamp 1663859327
transform 1 0 80304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_709
timestamp 1663859327
transform 1 0 80752 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_712
timestamp 1663859327
transform 1 0 81088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_776
timestamp 1663859327
transform 1 0 88256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_780
timestamp 1663859327
transform 1 0 88704 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_783
timestamp 1663859327
transform 1 0 89040 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_847
timestamp 1663859327
transform 1 0 96208 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_851
timestamp 1663859327
transform 1 0 96656 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_854
timestamp 1663859327
transform 1 0 96992 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_918
timestamp 1663859327
transform 1 0 104160 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_922
timestamp 1663859327
transform 1 0 104608 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_925
timestamp 1663859327
transform 1 0 104944 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_989
timestamp 1663859327
transform 1 0 112112 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_993
timestamp 1663859327
transform 1 0 112560 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_996
timestamp 1663859327
transform 1 0 112896 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_1028
timestamp 1663859327
transform 1 0 116480 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_1044
timestamp 1663859327
transform 1 0 118272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1663859327
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_7
timestamp 1663859327
transform 1 0 2128 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_23
timestamp 1663859327
transform 1 0 3920 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_31
timestamp 1663859327
transform 1 0 4816 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1663859327
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1663859327
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1663859327
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1663859327
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1663859327
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1663859327
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1663859327
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1663859327
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1663859327
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1663859327
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1663859327
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1663859327
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1663859327
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1663859327
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1663859327
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1663859327
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_456
timestamp 1663859327
transform 1 0 52416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1663859327
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_463
timestamp 1663859327
transform 1 0 53200 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_495
timestamp 1663859327
transform 1 0 56784 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_511
timestamp 1663859327
transform 1 0 58576 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_515
timestamp 1663859327
transform 1 0 59024 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_517
timestamp 1663859327
transform 1 0 59248 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_520
timestamp 1663859327
transform 1 0 59584 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_528
timestamp 1663859327
transform 1 0 60480 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_534
timestamp 1663859327
transform 1 0 61152 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_598
timestamp 1663859327
transform 1 0 68320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_602
timestamp 1663859327
transform 1 0 68768 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_605
timestamp 1663859327
transform 1 0 69104 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_669
timestamp 1663859327
transform 1 0 76272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_673
timestamp 1663859327
transform 1 0 76720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_676
timestamp 1663859327
transform 1 0 77056 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_740
timestamp 1663859327
transform 1 0 84224 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_744
timestamp 1663859327
transform 1 0 84672 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_747
timestamp 1663859327
transform 1 0 85008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_811
timestamp 1663859327
transform 1 0 92176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_815
timestamp 1663859327
transform 1 0 92624 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_818
timestamp 1663859327
transform 1 0 92960 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_882
timestamp 1663859327
transform 1 0 100128 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_886
timestamp 1663859327
transform 1 0 100576 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_889
timestamp 1663859327
transform 1 0 100912 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_953
timestamp 1663859327
transform 1 0 108080 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_957
timestamp 1663859327
transform 1 0 108528 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_960
timestamp 1663859327
transform 1 0 108864 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_1024
timestamp 1663859327
transform 1 0 116032 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1028
timestamp 1663859327
transform 1 0 116480 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_1031
timestamp 1663859327
transform 1 0 116816 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1039
timestamp 1663859327
transform 1 0 117712 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_1044
timestamp 1663859327
transform 1 0 118272 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_2
timestamp 1663859327
transform 1 0 1568 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_7
timestamp 1663859327
transform 1 0 2128 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1663859327
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1663859327
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1663859327
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1663859327
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1663859327
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1663859327
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1663859327
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1663859327
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1663859327
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1663859327
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1663859327
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1663859327
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_357
timestamp 1663859327
transform 1 0 41328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_421
timestamp 1663859327
transform 1 0 48496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1663859327
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1663859327
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_492
timestamp 1663859327
transform 1 0 56448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1663859327
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_499
timestamp 1663859327
transform 1 0 57232 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_563
timestamp 1663859327
transform 1 0 64400 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_567
timestamp 1663859327
transform 1 0 64848 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_570
timestamp 1663859327
transform 1 0 65184 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_634
timestamp 1663859327
transform 1 0 72352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_638
timestamp 1663859327
transform 1 0 72800 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_641
timestamp 1663859327
transform 1 0 73136 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_705
timestamp 1663859327
transform 1 0 80304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_709
timestamp 1663859327
transform 1 0 80752 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_712
timestamp 1663859327
transform 1 0 81088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_776
timestamp 1663859327
transform 1 0 88256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_780
timestamp 1663859327
transform 1 0 88704 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_783
timestamp 1663859327
transform 1 0 89040 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_847
timestamp 1663859327
transform 1 0 96208 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_851
timestamp 1663859327
transform 1 0 96656 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_854
timestamp 1663859327
transform 1 0 96992 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_918
timestamp 1663859327
transform 1 0 104160 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_922
timestamp 1663859327
transform 1 0 104608 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_925
timestamp 1663859327
transform 1 0 104944 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_989
timestamp 1663859327
transform 1 0 112112 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_993
timestamp 1663859327
transform 1 0 112560 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_996
timestamp 1663859327
transform 1 0 112896 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_1028
timestamp 1663859327
transform 1 0 116480 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_1044
timestamp 1663859327
transform 1 0 118272 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1663859327
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1663859327
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1663859327
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1663859327
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1663859327
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1663859327
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1663859327
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1663859327
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1663859327
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1663859327
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1663859327
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1663859327
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1663859327
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1663859327
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1663859327
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1663859327
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1663859327
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_392
timestamp 1663859327
transform 1 0 45248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_456
timestamp 1663859327
transform 1 0 52416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1663859327
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_463
timestamp 1663859327
transform 1 0 53200 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_527
timestamp 1663859327
transform 1 0 60368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_531
timestamp 1663859327
transform 1 0 60816 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_534
timestamp 1663859327
transform 1 0 61152 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_598
timestamp 1663859327
transform 1 0 68320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_602
timestamp 1663859327
transform 1 0 68768 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_605
timestamp 1663859327
transform 1 0 69104 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_669
timestamp 1663859327
transform 1 0 76272 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_673
timestamp 1663859327
transform 1 0 76720 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_676
timestamp 1663859327
transform 1 0 77056 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_740
timestamp 1663859327
transform 1 0 84224 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_744
timestamp 1663859327
transform 1 0 84672 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_747
timestamp 1663859327
transform 1 0 85008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_811
timestamp 1663859327
transform 1 0 92176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_815
timestamp 1663859327
transform 1 0 92624 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_818
timestamp 1663859327
transform 1 0 92960 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_882
timestamp 1663859327
transform 1 0 100128 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_886
timestamp 1663859327
transform 1 0 100576 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_889
timestamp 1663859327
transform 1 0 100912 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_953
timestamp 1663859327
transform 1 0 108080 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_957
timestamp 1663859327
transform 1 0 108528 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_960
timestamp 1663859327
transform 1 0 108864 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1024
timestamp 1663859327
transform 1 0 116032 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_1028
timestamp 1663859327
transform 1 0 116480 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_1031
timestamp 1663859327
transform 1 0 116816 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_1039
timestamp 1663859327
transform 1 0 117712 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_1043
timestamp 1663859327
transform 1 0 118160 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1663859327
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1663859327
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1663859327
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1663859327
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1663859327
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1663859327
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1663859327
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1663859327
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1663859327
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1663859327
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1663859327
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1663859327
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1663859327
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1663859327
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1663859327
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_357
timestamp 1663859327
transform 1 0 41328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_421
timestamp 1663859327
transform 1 0 48496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1663859327
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1663859327
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1663859327
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1663859327
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_499
timestamp 1663859327
transform 1 0 57232 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_563
timestamp 1663859327
transform 1 0 64400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_567
timestamp 1663859327
transform 1 0 64848 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_570
timestamp 1663859327
transform 1 0 65184 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_634
timestamp 1663859327
transform 1 0 72352 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_638
timestamp 1663859327
transform 1 0 72800 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_641
timestamp 1663859327
transform 1 0 73136 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_705
timestamp 1663859327
transform 1 0 80304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_709
timestamp 1663859327
transform 1 0 80752 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_712
timestamp 1663859327
transform 1 0 81088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_776
timestamp 1663859327
transform 1 0 88256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_780
timestamp 1663859327
transform 1 0 88704 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_783
timestamp 1663859327
transform 1 0 89040 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_847
timestamp 1663859327
transform 1 0 96208 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_851
timestamp 1663859327
transform 1 0 96656 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_854
timestamp 1663859327
transform 1 0 96992 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_918
timestamp 1663859327
transform 1 0 104160 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_922
timestamp 1663859327
transform 1 0 104608 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_925
timestamp 1663859327
transform 1 0 104944 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_989
timestamp 1663859327
transform 1 0 112112 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_993
timestamp 1663859327
transform 1 0 112560 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_996
timestamp 1663859327
transform 1 0 112896 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_1028
timestamp 1663859327
transform 1 0 116480 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_1044
timestamp 1663859327
transform 1 0 118272 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1663859327
transform 1 0 1568 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_5
timestamp 1663859327
transform 1 0 1904 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_21
timestamp 1663859327
transform 1 0 3696 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_29
timestamp 1663859327
transform 1 0 4592 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_33
timestamp 1663859327
transform 1 0 5040 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1663859327
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1663859327
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1663859327
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1663859327
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1663859327
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1663859327
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1663859327
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1663859327
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1663859327
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1663859327
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1663859327
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1663859327
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1663859327
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1663859327
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1663859327
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_392
timestamp 1663859327
transform 1 0 45248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_456
timestamp 1663859327
transform 1 0 52416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1663859327
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_463
timestamp 1663859327
transform 1 0 53200 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_527
timestamp 1663859327
transform 1 0 60368 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_531
timestamp 1663859327
transform 1 0 60816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_534
timestamp 1663859327
transform 1 0 61152 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_598
timestamp 1663859327
transform 1 0 68320 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_602
timestamp 1663859327
transform 1 0 68768 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_605
timestamp 1663859327
transform 1 0 69104 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_669
timestamp 1663859327
transform 1 0 76272 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_673
timestamp 1663859327
transform 1 0 76720 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_676
timestamp 1663859327
transform 1 0 77056 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_740
timestamp 1663859327
transform 1 0 84224 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_744
timestamp 1663859327
transform 1 0 84672 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_747
timestamp 1663859327
transform 1 0 85008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_811
timestamp 1663859327
transform 1 0 92176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_815
timestamp 1663859327
transform 1 0 92624 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_818
timestamp 1663859327
transform 1 0 92960 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_882
timestamp 1663859327
transform 1 0 100128 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_886
timestamp 1663859327
transform 1 0 100576 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_889
timestamp 1663859327
transform 1 0 100912 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_953
timestamp 1663859327
transform 1 0 108080 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_957
timestamp 1663859327
transform 1 0 108528 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_960
timestamp 1663859327
transform 1 0 108864 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_1024
timestamp 1663859327
transform 1 0 116032 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1028
timestamp 1663859327
transform 1 0 116480 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_1031
timestamp 1663859327
transform 1 0 116816 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1039
timestamp 1663859327
transform 1 0 117712 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_1044
timestamp 1663859327
transform 1 0 118272 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1663859327
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_9
timestamp 1663859327
transform 1 0 2352 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_41
timestamp 1663859327
transform 1 0 5936 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_57
timestamp 1663859327
transform 1 0 7728 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_65
timestamp 1663859327
transform 1 0 8624 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_69
timestamp 1663859327
transform 1 0 9072 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1663859327
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1663859327
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1663859327
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1663859327
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1663859327
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1663859327
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1663859327
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1663859327
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1663859327
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1663859327
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1663859327
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1663859327
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_357
timestamp 1663859327
transform 1 0 41328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_421
timestamp 1663859327
transform 1 0 48496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1663859327
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1663859327
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_492
timestamp 1663859327
transform 1 0 56448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1663859327
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_499
timestamp 1663859327
transform 1 0 57232 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_563
timestamp 1663859327
transform 1 0 64400 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_567
timestamp 1663859327
transform 1 0 64848 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_570
timestamp 1663859327
transform 1 0 65184 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_634
timestamp 1663859327
transform 1 0 72352 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_638
timestamp 1663859327
transform 1 0 72800 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_641
timestamp 1663859327
transform 1 0 73136 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_705
timestamp 1663859327
transform 1 0 80304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_709
timestamp 1663859327
transform 1 0 80752 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_712
timestamp 1663859327
transform 1 0 81088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_776
timestamp 1663859327
transform 1 0 88256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_780
timestamp 1663859327
transform 1 0 88704 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_783
timestamp 1663859327
transform 1 0 89040 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_847
timestamp 1663859327
transform 1 0 96208 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_851
timestamp 1663859327
transform 1 0 96656 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_854
timestamp 1663859327
transform 1 0 96992 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_918
timestamp 1663859327
transform 1 0 104160 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_922
timestamp 1663859327
transform 1 0 104608 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_925
timestamp 1663859327
transform 1 0 104944 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_989
timestamp 1663859327
transform 1 0 112112 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_993
timestamp 1663859327
transform 1 0 112560 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_996
timestamp 1663859327
transform 1 0 112896 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_1028
timestamp 1663859327
transform 1 0 116480 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_1044
timestamp 1663859327
transform 1 0 118272 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1663859327
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_9
timestamp 1663859327
transform 1 0 2352 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_13
timestamp 1663859327
transform 1 0 2800 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_29
timestamp 1663859327
transform 1 0 4592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_33
timestamp 1663859327
transform 1 0 5040 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1663859327
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1663859327
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1663859327
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1663859327
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1663859327
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1663859327
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1663859327
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1663859327
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1663859327
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1663859327
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1663859327
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1663859327
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1663859327
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1663859327
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1663859327
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_392
timestamp 1663859327
transform 1 0 45248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_456
timestamp 1663859327
transform 1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1663859327
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_463
timestamp 1663859327
transform 1 0 53200 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_527
timestamp 1663859327
transform 1 0 60368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_531
timestamp 1663859327
transform 1 0 60816 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_534
timestamp 1663859327
transform 1 0 61152 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_598
timestamp 1663859327
transform 1 0 68320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_602
timestamp 1663859327
transform 1 0 68768 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_605
timestamp 1663859327
transform 1 0 69104 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_669
timestamp 1663859327
transform 1 0 76272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_673
timestamp 1663859327
transform 1 0 76720 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_676
timestamp 1663859327
transform 1 0 77056 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_740
timestamp 1663859327
transform 1 0 84224 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_744
timestamp 1663859327
transform 1 0 84672 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_747
timestamp 1663859327
transform 1 0 85008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_811
timestamp 1663859327
transform 1 0 92176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_815
timestamp 1663859327
transform 1 0 92624 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_818
timestamp 1663859327
transform 1 0 92960 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_882
timestamp 1663859327
transform 1 0 100128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_886
timestamp 1663859327
transform 1 0 100576 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_889
timestamp 1663859327
transform 1 0 100912 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_953
timestamp 1663859327
transform 1 0 108080 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_957
timestamp 1663859327
transform 1 0 108528 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_960
timestamp 1663859327
transform 1 0 108864 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_1024
timestamp 1663859327
transform 1 0 116032 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1028
timestamp 1663859327
transform 1 0 116480 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_1031
timestamp 1663859327
transform 1 0 116816 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1039
timestamp 1663859327
transform 1 0 117712 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_1044
timestamp 1663859327
transform 1 0 118272 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_2
timestamp 1663859327
transform 1 0 1568 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_7
timestamp 1663859327
transform 1 0 2128 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1663859327
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1663859327
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1663859327
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1663859327
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1663859327
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1663859327
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1663859327
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1663859327
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1663859327
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1663859327
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1663859327
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1663859327
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_357
timestamp 1663859327
transform 1 0 41328 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_421
timestamp 1663859327
transform 1 0 48496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1663859327
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_428
timestamp 1663859327
transform 1 0 49280 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_492
timestamp 1663859327
transform 1 0 56448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1663859327
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_499
timestamp 1663859327
transform 1 0 57232 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_563
timestamp 1663859327
transform 1 0 64400 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_567
timestamp 1663859327
transform 1 0 64848 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_570
timestamp 1663859327
transform 1 0 65184 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_634
timestamp 1663859327
transform 1 0 72352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_638
timestamp 1663859327
transform 1 0 72800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_641
timestamp 1663859327
transform 1 0 73136 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_705
timestamp 1663859327
transform 1 0 80304 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_709
timestamp 1663859327
transform 1 0 80752 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_712
timestamp 1663859327
transform 1 0 81088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_776
timestamp 1663859327
transform 1 0 88256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_780
timestamp 1663859327
transform 1 0 88704 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_783
timestamp 1663859327
transform 1 0 89040 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_847
timestamp 1663859327
transform 1 0 96208 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_851
timestamp 1663859327
transform 1 0 96656 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_854
timestamp 1663859327
transform 1 0 96992 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_918
timestamp 1663859327
transform 1 0 104160 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_922
timestamp 1663859327
transform 1 0 104608 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_925
timestamp 1663859327
transform 1 0 104944 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_989
timestamp 1663859327
transform 1 0 112112 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_993
timestamp 1663859327
transform 1 0 112560 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_996
timestamp 1663859327
transform 1 0 112896 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_1028
timestamp 1663859327
transform 1 0 116480 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_1044
timestamp 1663859327
transform 1 0 118272 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1663859327
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1663859327
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1663859327
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1663859327
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1663859327
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1663859327
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1663859327
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1663859327
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1663859327
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1663859327
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1663859327
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1663859327
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1663859327
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1663859327
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1663859327
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1663859327
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1663859327
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_392
timestamp 1663859327
transform 1 0 45248 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_456
timestamp 1663859327
transform 1 0 52416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1663859327
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_463
timestamp 1663859327
transform 1 0 53200 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_527
timestamp 1663859327
transform 1 0 60368 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_531
timestamp 1663859327
transform 1 0 60816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_534
timestamp 1663859327
transform 1 0 61152 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_598
timestamp 1663859327
transform 1 0 68320 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_602
timestamp 1663859327
transform 1 0 68768 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_605
timestamp 1663859327
transform 1 0 69104 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_669
timestamp 1663859327
transform 1 0 76272 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_673
timestamp 1663859327
transform 1 0 76720 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_676
timestamp 1663859327
transform 1 0 77056 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_740
timestamp 1663859327
transform 1 0 84224 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_744
timestamp 1663859327
transform 1 0 84672 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_747
timestamp 1663859327
transform 1 0 85008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_811
timestamp 1663859327
transform 1 0 92176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_815
timestamp 1663859327
transform 1 0 92624 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_818
timestamp 1663859327
transform 1 0 92960 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_882
timestamp 1663859327
transform 1 0 100128 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_886
timestamp 1663859327
transform 1 0 100576 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_889
timestamp 1663859327
transform 1 0 100912 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_953
timestamp 1663859327
transform 1 0 108080 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_957
timestamp 1663859327
transform 1 0 108528 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_960
timestamp 1663859327
transform 1 0 108864 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_1024
timestamp 1663859327
transform 1 0 116032 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1028
timestamp 1663859327
transform 1 0 116480 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_1031
timestamp 1663859327
transform 1 0 116816 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1039
timestamp 1663859327
transform 1 0 117712 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_1044
timestamp 1663859327
transform 1 0 118272 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_2
timestamp 1663859327
transform 1 0 1568 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_17
timestamp 1663859327
transform 1 0 3248 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_21
timestamp 1663859327
transform 1 0 3696 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_53
timestamp 1663859327
transform 1 0 7280 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_69
timestamp 1663859327
transform 1 0 9072 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1663859327
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1663859327
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1663859327
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1663859327
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1663859327
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1663859327
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1663859327
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1663859327
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1663859327
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1663859327
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1663859327
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1663859327
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_357
timestamp 1663859327
transform 1 0 41328 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_421
timestamp 1663859327
transform 1 0 48496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1663859327
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_428
timestamp 1663859327
transform 1 0 49280 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_492
timestamp 1663859327
transform 1 0 56448 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1663859327
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_499
timestamp 1663859327
transform 1 0 57232 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_563
timestamp 1663859327
transform 1 0 64400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_567
timestamp 1663859327
transform 1 0 64848 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_570
timestamp 1663859327
transform 1 0 65184 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_634
timestamp 1663859327
transform 1 0 72352 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_638
timestamp 1663859327
transform 1 0 72800 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_641
timestamp 1663859327
transform 1 0 73136 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_705
timestamp 1663859327
transform 1 0 80304 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_709
timestamp 1663859327
transform 1 0 80752 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_712
timestamp 1663859327
transform 1 0 81088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_776
timestamp 1663859327
transform 1 0 88256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_780
timestamp 1663859327
transform 1 0 88704 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_783
timestamp 1663859327
transform 1 0 89040 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_847
timestamp 1663859327
transform 1 0 96208 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_851
timestamp 1663859327
transform 1 0 96656 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_854
timestamp 1663859327
transform 1 0 96992 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_918
timestamp 1663859327
transform 1 0 104160 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_922
timestamp 1663859327
transform 1 0 104608 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_925
timestamp 1663859327
transform 1 0 104944 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_989
timestamp 1663859327
transform 1 0 112112 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_993
timestamp 1663859327
transform 1 0 112560 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_996
timestamp 1663859327
transform 1 0 112896 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_1028
timestamp 1663859327
transform 1 0 116480 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_1044
timestamp 1663859327
transform 1 0 118272 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1663859327
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1663859327
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1663859327
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1663859327
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1663859327
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1663859327
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1663859327
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1663859327
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1663859327
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1663859327
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1663859327
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1663859327
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1663859327
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1663859327
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1663859327
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1663859327
transform 1 0 44464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1663859327
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_392
timestamp 1663859327
transform 1 0 45248 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_456
timestamp 1663859327
transform 1 0 52416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1663859327
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_463
timestamp 1663859327
transform 1 0 53200 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_527
timestamp 1663859327
transform 1 0 60368 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_531
timestamp 1663859327
transform 1 0 60816 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_534
timestamp 1663859327
transform 1 0 61152 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_598
timestamp 1663859327
transform 1 0 68320 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_602
timestamp 1663859327
transform 1 0 68768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_605
timestamp 1663859327
transform 1 0 69104 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_669
timestamp 1663859327
transform 1 0 76272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_673
timestamp 1663859327
transform 1 0 76720 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_676
timestamp 1663859327
transform 1 0 77056 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_740
timestamp 1663859327
transform 1 0 84224 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_744
timestamp 1663859327
transform 1 0 84672 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_747
timestamp 1663859327
transform 1 0 85008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_811
timestamp 1663859327
transform 1 0 92176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_815
timestamp 1663859327
transform 1 0 92624 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_818
timestamp 1663859327
transform 1 0 92960 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_882
timestamp 1663859327
transform 1 0 100128 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_886
timestamp 1663859327
transform 1 0 100576 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_889
timestamp 1663859327
transform 1 0 100912 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_953
timestamp 1663859327
transform 1 0 108080 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_957
timestamp 1663859327
transform 1 0 108528 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_960
timestamp 1663859327
transform 1 0 108864 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1024
timestamp 1663859327
transform 1 0 116032 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_1028
timestamp 1663859327
transform 1 0 116480 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_1031
timestamp 1663859327
transform 1 0 116816 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_1039
timestamp 1663859327
transform 1 0 117712 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_1043
timestamp 1663859327
transform 1 0 118160 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_2
timestamp 1663859327
transform 1 0 1568 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_7
timestamp 1663859327
transform 1 0 2128 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1663859327
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1663859327
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1663859327
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1663859327
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1663859327
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1663859327
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1663859327
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1663859327
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1663859327
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1663859327
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1663859327
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1663859327
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_357
timestamp 1663859327
transform 1 0 41328 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_421
timestamp 1663859327
transform 1 0 48496 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1663859327
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_428
timestamp 1663859327
transform 1 0 49280 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_492
timestamp 1663859327
transform 1 0 56448 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1663859327
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_499
timestamp 1663859327
transform 1 0 57232 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_563
timestamp 1663859327
transform 1 0 64400 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_567
timestamp 1663859327
transform 1 0 64848 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_570
timestamp 1663859327
transform 1 0 65184 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_634
timestamp 1663859327
transform 1 0 72352 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_638
timestamp 1663859327
transform 1 0 72800 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_641
timestamp 1663859327
transform 1 0 73136 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_705
timestamp 1663859327
transform 1 0 80304 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_709
timestamp 1663859327
transform 1 0 80752 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_712
timestamp 1663859327
transform 1 0 81088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_776
timestamp 1663859327
transform 1 0 88256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_780
timestamp 1663859327
transform 1 0 88704 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_783
timestamp 1663859327
transform 1 0 89040 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_847
timestamp 1663859327
transform 1 0 96208 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_851
timestamp 1663859327
transform 1 0 96656 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_854
timestamp 1663859327
transform 1 0 96992 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_918
timestamp 1663859327
transform 1 0 104160 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_922
timestamp 1663859327
transform 1 0 104608 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_925
timestamp 1663859327
transform 1 0 104944 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_989
timestamp 1663859327
transform 1 0 112112 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_993
timestamp 1663859327
transform 1 0 112560 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_996
timestamp 1663859327
transform 1 0 112896 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_1028
timestamp 1663859327
transform 1 0 116480 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_1044
timestamp 1663859327
transform 1 0 118272 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1663859327
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1663859327
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1663859327
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1663859327
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1663859327
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1663859327
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1663859327
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1663859327
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1663859327
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1663859327
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1663859327
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1663859327
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1663859327
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1663859327
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1663859327
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_385
timestamp 1663859327
transform 1 0 44464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1663859327
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_392
timestamp 1663859327
transform 1 0 45248 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_456
timestamp 1663859327
transform 1 0 52416 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1663859327
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_463
timestamp 1663859327
transform 1 0 53200 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_527
timestamp 1663859327
transform 1 0 60368 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_531
timestamp 1663859327
transform 1 0 60816 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_534
timestamp 1663859327
transform 1 0 61152 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_598
timestamp 1663859327
transform 1 0 68320 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_602
timestamp 1663859327
transform 1 0 68768 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_605
timestamp 1663859327
transform 1 0 69104 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_669
timestamp 1663859327
transform 1 0 76272 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_673
timestamp 1663859327
transform 1 0 76720 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_676
timestamp 1663859327
transform 1 0 77056 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_740
timestamp 1663859327
transform 1 0 84224 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_744
timestamp 1663859327
transform 1 0 84672 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_747
timestamp 1663859327
transform 1 0 85008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_811
timestamp 1663859327
transform 1 0 92176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_815
timestamp 1663859327
transform 1 0 92624 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_818
timestamp 1663859327
transform 1 0 92960 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_882
timestamp 1663859327
transform 1 0 100128 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_886
timestamp 1663859327
transform 1 0 100576 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_889
timestamp 1663859327
transform 1 0 100912 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_953
timestamp 1663859327
transform 1 0 108080 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_957
timestamp 1663859327
transform 1 0 108528 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_960
timestamp 1663859327
transform 1 0 108864 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1024
timestamp 1663859327
transform 1 0 116032 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_1028
timestamp 1663859327
transform 1 0 116480 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_1031
timestamp 1663859327
transform 1 0 116816 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_1039
timestamp 1663859327
transform 1 0 117712 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_1043
timestamp 1663859327
transform 1 0 118160 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1663859327
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1663859327
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1663859327
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1663859327
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1663859327
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1663859327
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1663859327
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1663859327
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1663859327
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1663859327
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1663859327
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1663859327
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1663859327
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1663859327
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1663859327
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_357
timestamp 1663859327
transform 1 0 41328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_421
timestamp 1663859327
transform 1 0 48496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1663859327
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_428
timestamp 1663859327
transform 1 0 49280 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_492
timestamp 1663859327
transform 1 0 56448 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1663859327
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_499
timestamp 1663859327
transform 1 0 57232 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_563
timestamp 1663859327
transform 1 0 64400 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_567
timestamp 1663859327
transform 1 0 64848 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_570
timestamp 1663859327
transform 1 0 65184 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_634
timestamp 1663859327
transform 1 0 72352 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_638
timestamp 1663859327
transform 1 0 72800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_641
timestamp 1663859327
transform 1 0 73136 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_705
timestamp 1663859327
transform 1 0 80304 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_709
timestamp 1663859327
transform 1 0 80752 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_712
timestamp 1663859327
transform 1 0 81088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_776
timestamp 1663859327
transform 1 0 88256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_780
timestamp 1663859327
transform 1 0 88704 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_783
timestamp 1663859327
transform 1 0 89040 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_847
timestamp 1663859327
transform 1 0 96208 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_851
timestamp 1663859327
transform 1 0 96656 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_854
timestamp 1663859327
transform 1 0 96992 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_918
timestamp 1663859327
transform 1 0 104160 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_922
timestamp 1663859327
transform 1 0 104608 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_925
timestamp 1663859327
transform 1 0 104944 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_989
timestamp 1663859327
transform 1 0 112112 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_993
timestamp 1663859327
transform 1 0 112560 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_996
timestamp 1663859327
transform 1 0 112896 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_1028
timestamp 1663859327
transform 1 0 116480 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_1044
timestamp 1663859327
transform 1 0 118272 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_2
timestamp 1663859327
transform 1 0 1568 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_5
timestamp 1663859327
transform 1 0 1904 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_21
timestamp 1663859327
transform 1 0 3696 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_29
timestamp 1663859327
transform 1 0 4592 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_33
timestamp 1663859327
transform 1 0 5040 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1663859327
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1663859327
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1663859327
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1663859327
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1663859327
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1663859327
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1663859327
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1663859327
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1663859327
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1663859327
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1663859327
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1663859327
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1663859327
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1663859327
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1663859327
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_392
timestamp 1663859327
transform 1 0 45248 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_456
timestamp 1663859327
transform 1 0 52416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1663859327
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_463
timestamp 1663859327
transform 1 0 53200 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_527
timestamp 1663859327
transform 1 0 60368 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_531
timestamp 1663859327
transform 1 0 60816 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_534
timestamp 1663859327
transform 1 0 61152 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_598
timestamp 1663859327
transform 1 0 68320 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_602
timestamp 1663859327
transform 1 0 68768 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_605
timestamp 1663859327
transform 1 0 69104 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_669
timestamp 1663859327
transform 1 0 76272 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_673
timestamp 1663859327
transform 1 0 76720 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_676
timestamp 1663859327
transform 1 0 77056 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_740
timestamp 1663859327
transform 1 0 84224 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_744
timestamp 1663859327
transform 1 0 84672 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_747
timestamp 1663859327
transform 1 0 85008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_811
timestamp 1663859327
transform 1 0 92176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_815
timestamp 1663859327
transform 1 0 92624 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_818
timestamp 1663859327
transform 1 0 92960 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_882
timestamp 1663859327
transform 1 0 100128 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_886
timestamp 1663859327
transform 1 0 100576 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_889
timestamp 1663859327
transform 1 0 100912 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_953
timestamp 1663859327
transform 1 0 108080 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_957
timestamp 1663859327
transform 1 0 108528 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_960
timestamp 1663859327
transform 1 0 108864 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1024
timestamp 1663859327
transform 1 0 116032 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_1028
timestamp 1663859327
transform 1 0 116480 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_1031
timestamp 1663859327
transform 1 0 116816 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_1039
timestamp 1663859327
transform 1 0 117712 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_1043
timestamp 1663859327
transform 1 0 118160 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_2
timestamp 1663859327
transform 1 0 1568 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_9
timestamp 1663859327
transform 1 0 2352 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_41
timestamp 1663859327
transform 1 0 5936 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_57
timestamp 1663859327
transform 1 0 7728 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_65
timestamp 1663859327
transform 1 0 8624 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_69
timestamp 1663859327
transform 1 0 9072 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1663859327
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1663859327
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1663859327
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1663859327
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1663859327
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1663859327
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1663859327
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1663859327
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1663859327
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1663859327
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1663859327
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1663859327
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_357
timestamp 1663859327
transform 1 0 41328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_421
timestamp 1663859327
transform 1 0 48496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1663859327
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1663859327
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_492
timestamp 1663859327
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1663859327
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_499
timestamp 1663859327
transform 1 0 57232 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_563
timestamp 1663859327
transform 1 0 64400 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_567
timestamp 1663859327
transform 1 0 64848 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_570
timestamp 1663859327
transform 1 0 65184 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_634
timestamp 1663859327
transform 1 0 72352 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_638
timestamp 1663859327
transform 1 0 72800 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_641
timestamp 1663859327
transform 1 0 73136 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_705
timestamp 1663859327
transform 1 0 80304 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_709
timestamp 1663859327
transform 1 0 80752 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_712
timestamp 1663859327
transform 1 0 81088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_776
timestamp 1663859327
transform 1 0 88256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_780
timestamp 1663859327
transform 1 0 88704 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_783
timestamp 1663859327
transform 1 0 89040 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_847
timestamp 1663859327
transform 1 0 96208 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_851
timestamp 1663859327
transform 1 0 96656 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_854
timestamp 1663859327
transform 1 0 96992 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_918
timestamp 1663859327
transform 1 0 104160 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_922
timestamp 1663859327
transform 1 0 104608 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_925
timestamp 1663859327
transform 1 0 104944 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_989
timestamp 1663859327
transform 1 0 112112 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_993
timestamp 1663859327
transform 1 0 112560 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_996
timestamp 1663859327
transform 1 0 112896 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_1028
timestamp 1663859327
transform 1 0 116480 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_1036
timestamp 1663859327
transform 1 0 117376 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_1044
timestamp 1663859327
transform 1 0 118272 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1663859327
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1663859327
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1663859327
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1663859327
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1663859327
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1663859327
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1663859327
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1663859327
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1663859327
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1663859327
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1663859327
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1663859327
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1663859327
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1663859327
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1663859327
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1663859327
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1663859327
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_392
timestamp 1663859327
transform 1 0 45248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_456
timestamp 1663859327
transform 1 0 52416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1663859327
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_463
timestamp 1663859327
transform 1 0 53200 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_527
timestamp 1663859327
transform 1 0 60368 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_531
timestamp 1663859327
transform 1 0 60816 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_534
timestamp 1663859327
transform 1 0 61152 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_598
timestamp 1663859327
transform 1 0 68320 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_602
timestamp 1663859327
transform 1 0 68768 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_605
timestamp 1663859327
transform 1 0 69104 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_669
timestamp 1663859327
transform 1 0 76272 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_673
timestamp 1663859327
transform 1 0 76720 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_676
timestamp 1663859327
transform 1 0 77056 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_740
timestamp 1663859327
transform 1 0 84224 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_744
timestamp 1663859327
transform 1 0 84672 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_747
timestamp 1663859327
transform 1 0 85008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_811
timestamp 1663859327
transform 1 0 92176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_815
timestamp 1663859327
transform 1 0 92624 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_818
timestamp 1663859327
transform 1 0 92960 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_882
timestamp 1663859327
transform 1 0 100128 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_886
timestamp 1663859327
transform 1 0 100576 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_889
timestamp 1663859327
transform 1 0 100912 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_953
timestamp 1663859327
transform 1 0 108080 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_957
timestamp 1663859327
transform 1 0 108528 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_960
timestamp 1663859327
transform 1 0 108864 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_1024
timestamp 1663859327
transform 1 0 116032 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1028
timestamp 1663859327
transform 1 0 116480 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_1031
timestamp 1663859327
transform 1 0 116816 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1039
timestamp 1663859327
transform 1 0 117712 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_1044
timestamp 1663859327
transform 1 0 118272 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1663859327
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1663859327
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1663859327
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1663859327
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1663859327
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1663859327
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1663859327
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1663859327
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1663859327
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1663859327
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1663859327
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1663859327
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1663859327
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1663859327
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1663859327
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1663859327
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_421
timestamp 1663859327
transform 1 0 48496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1663859327
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1663859327
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_492
timestamp 1663859327
transform 1 0 56448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1663859327
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_499
timestamp 1663859327
transform 1 0 57232 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_563
timestamp 1663859327
transform 1 0 64400 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_567
timestamp 1663859327
transform 1 0 64848 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_570
timestamp 1663859327
transform 1 0 65184 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_634
timestamp 1663859327
transform 1 0 72352 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_638
timestamp 1663859327
transform 1 0 72800 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_641
timestamp 1663859327
transform 1 0 73136 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_705
timestamp 1663859327
transform 1 0 80304 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_709
timestamp 1663859327
transform 1 0 80752 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_712
timestamp 1663859327
transform 1 0 81088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_776
timestamp 1663859327
transform 1 0 88256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_780
timestamp 1663859327
transform 1 0 88704 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_783
timestamp 1663859327
transform 1 0 89040 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_847
timestamp 1663859327
transform 1 0 96208 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_851
timestamp 1663859327
transform 1 0 96656 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_854
timestamp 1663859327
transform 1 0 96992 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_918
timestamp 1663859327
transform 1 0 104160 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_922
timestamp 1663859327
transform 1 0 104608 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_925
timestamp 1663859327
transform 1 0 104944 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_989
timestamp 1663859327
transform 1 0 112112 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_993
timestamp 1663859327
transform 1 0 112560 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_996
timestamp 1663859327
transform 1 0 112896 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_1028
timestamp 1663859327
transform 1 0 116480 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_1044
timestamp 1663859327
transform 1 0 118272 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1663859327
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1663859327
transform 1 0 5152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1663859327
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1663859327
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1663859327
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1663859327
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1663859327
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1663859327
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1663859327
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1663859327
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1663859327
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1663859327
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1663859327
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1663859327
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1663859327
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1663859327
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1663859327
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_392
timestamp 1663859327
transform 1 0 45248 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_456
timestamp 1663859327
transform 1 0 52416 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1663859327
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_463
timestamp 1663859327
transform 1 0 53200 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_527
timestamp 1663859327
transform 1 0 60368 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_531
timestamp 1663859327
transform 1 0 60816 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_534
timestamp 1663859327
transform 1 0 61152 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_598
timestamp 1663859327
transform 1 0 68320 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_602
timestamp 1663859327
transform 1 0 68768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_605
timestamp 1663859327
transform 1 0 69104 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_669
timestamp 1663859327
transform 1 0 76272 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_673
timestamp 1663859327
transform 1 0 76720 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_676
timestamp 1663859327
transform 1 0 77056 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_740
timestamp 1663859327
transform 1 0 84224 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_744
timestamp 1663859327
transform 1 0 84672 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_747
timestamp 1663859327
transform 1 0 85008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_811
timestamp 1663859327
transform 1 0 92176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_815
timestamp 1663859327
transform 1 0 92624 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_818
timestamp 1663859327
transform 1 0 92960 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_882
timestamp 1663859327
transform 1 0 100128 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_886
timestamp 1663859327
transform 1 0 100576 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_889
timestamp 1663859327
transform 1 0 100912 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_953
timestamp 1663859327
transform 1 0 108080 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_957
timestamp 1663859327
transform 1 0 108528 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_960
timestamp 1663859327
transform 1 0 108864 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1024
timestamp 1663859327
transform 1 0 116032 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_1028
timestamp 1663859327
transform 1 0 116480 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_1031
timestamp 1663859327
transform 1 0 116816 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_1039
timestamp 1663859327
transform 1 0 117712 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_1043
timestamp 1663859327
transform 1 0 118160 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1663859327
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1663859327
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_70
timestamp 1663859327
transform 1 0 9184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_73
timestamp 1663859327
transform 1 0 9520 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_137
timestamp 1663859327
transform 1 0 16688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1663859327
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1663859327
transform 1 0 17472 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_208
timestamp 1663859327
transform 1 0 24640 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1663859327
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1663859327
transform 1 0 25424 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_279
timestamp 1663859327
transform 1 0 32592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1663859327
transform 1 0 33040 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1663859327
transform 1 0 33376 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1663859327
transform 1 0 40544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1663859327
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_357
timestamp 1663859327
transform 1 0 41328 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_421
timestamp 1663859327
transform 1 0 48496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_425
timestamp 1663859327
transform 1 0 48944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_428
timestamp 1663859327
transform 1 0 49280 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_492
timestamp 1663859327
transform 1 0 56448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1663859327
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_499
timestamp 1663859327
transform 1 0 57232 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_563
timestamp 1663859327
transform 1 0 64400 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_567
timestamp 1663859327
transform 1 0 64848 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_570
timestamp 1663859327
transform 1 0 65184 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_634
timestamp 1663859327
transform 1 0 72352 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_638
timestamp 1663859327
transform 1 0 72800 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_641
timestamp 1663859327
transform 1 0 73136 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_705
timestamp 1663859327
transform 1 0 80304 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_709
timestamp 1663859327
transform 1 0 80752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_712
timestamp 1663859327
transform 1 0 81088 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_776
timestamp 1663859327
transform 1 0 88256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_780
timestamp 1663859327
transform 1 0 88704 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_783
timestamp 1663859327
transform 1 0 89040 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_847
timestamp 1663859327
transform 1 0 96208 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_851
timestamp 1663859327
transform 1 0 96656 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_854
timestamp 1663859327
transform 1 0 96992 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_918
timestamp 1663859327
transform 1 0 104160 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_922
timestamp 1663859327
transform 1 0 104608 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_925
timestamp 1663859327
transform 1 0 104944 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_989
timestamp 1663859327
transform 1 0 112112 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_993
timestamp 1663859327
transform 1 0 112560 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_996
timestamp 1663859327
transform 1 0 112896 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_1028
timestamp 1663859327
transform 1 0 116480 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_1044
timestamp 1663859327
transform 1 0 118272 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_2
timestamp 1663859327
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1663859327
transform 1 0 5152 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1663859327
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1663859327
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1663859327
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_108
timestamp 1663859327
transform 1 0 13440 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_172
timestamp 1663859327
transform 1 0 20608 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1663859327
transform 1 0 21056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1663859327
transform 1 0 21392 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_243
timestamp 1663859327
transform 1 0 28560 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1663859327
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1663859327
transform 1 0 29344 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_314
timestamp 1663859327
transform 1 0 36512 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1663859327
transform 1 0 36960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_321
timestamp 1663859327
transform 1 0 37296 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_385
timestamp 1663859327
transform 1 0 44464 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1663859327
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_392
timestamp 1663859327
transform 1 0 45248 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_456
timestamp 1663859327
transform 1 0 52416 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1663859327
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_463
timestamp 1663859327
transform 1 0 53200 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_527
timestamp 1663859327
transform 1 0 60368 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_531
timestamp 1663859327
transform 1 0 60816 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_534
timestamp 1663859327
transform 1 0 61152 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_598
timestamp 1663859327
transform 1 0 68320 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_602
timestamp 1663859327
transform 1 0 68768 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_605
timestamp 1663859327
transform 1 0 69104 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_669
timestamp 1663859327
transform 1 0 76272 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_673
timestamp 1663859327
transform 1 0 76720 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_676
timestamp 1663859327
transform 1 0 77056 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_740
timestamp 1663859327
transform 1 0 84224 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_744
timestamp 1663859327
transform 1 0 84672 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_747
timestamp 1663859327
transform 1 0 85008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_811
timestamp 1663859327
transform 1 0 92176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_815
timestamp 1663859327
transform 1 0 92624 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_818
timestamp 1663859327
transform 1 0 92960 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_882
timestamp 1663859327
transform 1 0 100128 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_886
timestamp 1663859327
transform 1 0 100576 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_889
timestamp 1663859327
transform 1 0 100912 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_953
timestamp 1663859327
transform 1 0 108080 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_957
timestamp 1663859327
transform 1 0 108528 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_960
timestamp 1663859327
transform 1 0 108864 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1024
timestamp 1663859327
transform 1 0 116032 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_1028
timestamp 1663859327
transform 1 0 116480 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_1031
timestamp 1663859327
transform 1 0 116816 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_1039
timestamp 1663859327
transform 1 0 117712 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_1043
timestamp 1663859327
transform 1 0 118160 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_2
timestamp 1663859327
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_66
timestamp 1663859327
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_70
timestamp 1663859327
transform 1 0 9184 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_73
timestamp 1663859327
transform 1 0 9520 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_137
timestamp 1663859327
transform 1 0 16688 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_141
timestamp 1663859327
transform 1 0 17136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1663859327
transform 1 0 17472 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_208
timestamp 1663859327
transform 1 0 24640 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1663859327
transform 1 0 25088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1663859327
transform 1 0 25424 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_279
timestamp 1663859327
transform 1 0 32592 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1663859327
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1663859327
transform 1 0 33376 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_350
timestamp 1663859327
transform 1 0 40544 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1663859327
transform 1 0 40992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_357
timestamp 1663859327
transform 1 0 41328 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_421
timestamp 1663859327
transform 1 0 48496 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_425
timestamp 1663859327
transform 1 0 48944 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_428
timestamp 1663859327
transform 1 0 49280 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_492
timestamp 1663859327
transform 1 0 56448 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_496
timestamp 1663859327
transform 1 0 56896 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_499
timestamp 1663859327
transform 1 0 57232 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_563
timestamp 1663859327
transform 1 0 64400 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_567
timestamp 1663859327
transform 1 0 64848 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_570
timestamp 1663859327
transform 1 0 65184 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_634
timestamp 1663859327
transform 1 0 72352 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_638
timestamp 1663859327
transform 1 0 72800 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_641
timestamp 1663859327
transform 1 0 73136 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_705
timestamp 1663859327
transform 1 0 80304 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_709
timestamp 1663859327
transform 1 0 80752 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_712
timestamp 1663859327
transform 1 0 81088 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_776
timestamp 1663859327
transform 1 0 88256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_780
timestamp 1663859327
transform 1 0 88704 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_783
timestamp 1663859327
transform 1 0 89040 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_847
timestamp 1663859327
transform 1 0 96208 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_851
timestamp 1663859327
transform 1 0 96656 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_854
timestamp 1663859327
transform 1 0 96992 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_918
timestamp 1663859327
transform 1 0 104160 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_922
timestamp 1663859327
transform 1 0 104608 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_925
timestamp 1663859327
transform 1 0 104944 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_989
timestamp 1663859327
transform 1 0 112112 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_993
timestamp 1663859327
transform 1 0 112560 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_996
timestamp 1663859327
transform 1 0 112896 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_1028
timestamp 1663859327
transform 1 0 116480 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_1036
timestamp 1663859327
transform 1 0 117376 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_1044
timestamp 1663859327
transform 1 0 118272 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_2
timestamp 1663859327
transform 1 0 1568 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_7
timestamp 1663859327
transform 1 0 2128 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_23
timestamp 1663859327
transform 1 0 3920 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_31
timestamp 1663859327
transform 1 0 4816 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_37
timestamp 1663859327
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_101
timestamp 1663859327
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1663859327
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_108
timestamp 1663859327
transform 1 0 13440 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_172
timestamp 1663859327
transform 1 0 20608 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1663859327
transform 1 0 21056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1663859327
transform 1 0 21392 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_243
timestamp 1663859327
transform 1 0 28560 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1663859327
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1663859327
transform 1 0 29344 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_314
timestamp 1663859327
transform 1 0 36512 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1663859327
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1663859327
transform 1 0 37296 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_385
timestamp 1663859327
transform 1 0 44464 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1663859327
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_392
timestamp 1663859327
transform 1 0 45248 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_456
timestamp 1663859327
transform 1 0 52416 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1663859327
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_463
timestamp 1663859327
transform 1 0 53200 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_527
timestamp 1663859327
transform 1 0 60368 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_531
timestamp 1663859327
transform 1 0 60816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_534
timestamp 1663859327
transform 1 0 61152 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_598
timestamp 1663859327
transform 1 0 68320 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_602
timestamp 1663859327
transform 1 0 68768 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_605
timestamp 1663859327
transform 1 0 69104 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_669
timestamp 1663859327
transform 1 0 76272 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_673
timestamp 1663859327
transform 1 0 76720 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_676
timestamp 1663859327
transform 1 0 77056 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_740
timestamp 1663859327
transform 1 0 84224 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_744
timestamp 1663859327
transform 1 0 84672 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_747
timestamp 1663859327
transform 1 0 85008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_811
timestamp 1663859327
transform 1 0 92176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_815
timestamp 1663859327
transform 1 0 92624 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_818
timestamp 1663859327
transform 1 0 92960 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_882
timestamp 1663859327
transform 1 0 100128 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_886
timestamp 1663859327
transform 1 0 100576 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_889
timestamp 1663859327
transform 1 0 100912 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_953
timestamp 1663859327
transform 1 0 108080 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_957
timestamp 1663859327
transform 1 0 108528 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_960
timestamp 1663859327
transform 1 0 108864 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1024
timestamp 1663859327
transform 1 0 116032 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_1028
timestamp 1663859327
transform 1 0 116480 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_1031
timestamp 1663859327
transform 1 0 116816 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_1039
timestamp 1663859327
transform 1 0 117712 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_1043
timestamp 1663859327
transform 1 0 118160 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_2
timestamp 1663859327
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_66
timestamp 1663859327
transform 1 0 8736 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_70
timestamp 1663859327
transform 1 0 9184 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_73
timestamp 1663859327
transform 1 0 9520 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_137
timestamp 1663859327
transform 1 0 16688 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1663859327
transform 1 0 17136 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_144
timestamp 1663859327
transform 1 0 17472 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_208
timestamp 1663859327
transform 1 0 24640 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1663859327
transform 1 0 25088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1663859327
transform 1 0 25424 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_279
timestamp 1663859327
transform 1 0 32592 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1663859327
transform 1 0 33040 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1663859327
transform 1 0 33376 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_350
timestamp 1663859327
transform 1 0 40544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1663859327
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_357
timestamp 1663859327
transform 1 0 41328 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_421
timestamp 1663859327
transform 1 0 48496 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_425
timestamp 1663859327
transform 1 0 48944 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_428
timestamp 1663859327
transform 1 0 49280 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_492
timestamp 1663859327
transform 1 0 56448 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_496
timestamp 1663859327
transform 1 0 56896 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_499
timestamp 1663859327
transform 1 0 57232 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_563
timestamp 1663859327
transform 1 0 64400 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_567
timestamp 1663859327
transform 1 0 64848 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_570
timestamp 1663859327
transform 1 0 65184 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_634
timestamp 1663859327
transform 1 0 72352 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_638
timestamp 1663859327
transform 1 0 72800 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_641
timestamp 1663859327
transform 1 0 73136 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_705
timestamp 1663859327
transform 1 0 80304 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_709
timestamp 1663859327
transform 1 0 80752 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_712
timestamp 1663859327
transform 1 0 81088 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_776
timestamp 1663859327
transform 1 0 88256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_780
timestamp 1663859327
transform 1 0 88704 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_783
timestamp 1663859327
transform 1 0 89040 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_847
timestamp 1663859327
transform 1 0 96208 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_851
timestamp 1663859327
transform 1 0 96656 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_854
timestamp 1663859327
transform 1 0 96992 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_918
timestamp 1663859327
transform 1 0 104160 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_922
timestamp 1663859327
transform 1 0 104608 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_925
timestamp 1663859327
transform 1 0 104944 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_989
timestamp 1663859327
transform 1 0 112112 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_993
timestamp 1663859327
transform 1 0 112560 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_996
timestamp 1663859327
transform 1 0 112896 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_1028
timestamp 1663859327
transform 1 0 116480 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_1036
timestamp 1663859327
transform 1 0 117376 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_1044
timestamp 1663859327
transform 1 0 118272 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_2
timestamp 1663859327
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_34
timestamp 1663859327
transform 1 0 5152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_37
timestamp 1663859327
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_101
timestamp 1663859327
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1663859327
transform 1 0 13104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_108
timestamp 1663859327
transform 1 0 13440 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_172
timestamp 1663859327
transform 1 0 20608 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1663859327
transform 1 0 21056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_179
timestamp 1663859327
transform 1 0 21392 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_243
timestamp 1663859327
transform 1 0 28560 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1663859327
transform 1 0 29008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1663859327
transform 1 0 29344 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_314
timestamp 1663859327
transform 1 0 36512 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1663859327
transform 1 0 36960 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1663859327
transform 1 0 37296 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_385
timestamp 1663859327
transform 1 0 44464 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1663859327
transform 1 0 44912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_392
timestamp 1663859327
transform 1 0 45248 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_456
timestamp 1663859327
transform 1 0 52416 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_460
timestamp 1663859327
transform 1 0 52864 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_463
timestamp 1663859327
transform 1 0 53200 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_527
timestamp 1663859327
transform 1 0 60368 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_531
timestamp 1663859327
transform 1 0 60816 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_534
timestamp 1663859327
transform 1 0 61152 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_598
timestamp 1663859327
transform 1 0 68320 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_602
timestamp 1663859327
transform 1 0 68768 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_605
timestamp 1663859327
transform 1 0 69104 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_669
timestamp 1663859327
transform 1 0 76272 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_673
timestamp 1663859327
transform 1 0 76720 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_676
timestamp 1663859327
transform 1 0 77056 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_740
timestamp 1663859327
transform 1 0 84224 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_744
timestamp 1663859327
transform 1 0 84672 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_747
timestamp 1663859327
transform 1 0 85008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_811
timestamp 1663859327
transform 1 0 92176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_815
timestamp 1663859327
transform 1 0 92624 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_818
timestamp 1663859327
transform 1 0 92960 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_882
timestamp 1663859327
transform 1 0 100128 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_886
timestamp 1663859327
transform 1 0 100576 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_889
timestamp 1663859327
transform 1 0 100912 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_953
timestamp 1663859327
transform 1 0 108080 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_957
timestamp 1663859327
transform 1 0 108528 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_960
timestamp 1663859327
transform 1 0 108864 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_1024
timestamp 1663859327
transform 1 0 116032 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1028
timestamp 1663859327
transform 1 0 116480 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_1031
timestamp 1663859327
transform 1 0 116816 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1039
timestamp 1663859327
transform 1 0 117712 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_1044
timestamp 1663859327
transform 1 0 118272 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_2
timestamp 1663859327
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_66
timestamp 1663859327
transform 1 0 8736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_70
timestamp 1663859327
transform 1 0 9184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_73
timestamp 1663859327
transform 1 0 9520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_137
timestamp 1663859327
transform 1 0 16688 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1663859327
transform 1 0 17136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_144
timestamp 1663859327
transform 1 0 17472 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_208
timestamp 1663859327
transform 1 0 24640 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_212
timestamp 1663859327
transform 1 0 25088 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_215
timestamp 1663859327
transform 1 0 25424 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_279
timestamp 1663859327
transform 1 0 32592 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_283
timestamp 1663859327
transform 1 0 33040 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1663859327
transform 1 0 33376 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_350
timestamp 1663859327
transform 1 0 40544 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1663859327
transform 1 0 40992 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_357
timestamp 1663859327
transform 1 0 41328 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_421
timestamp 1663859327
transform 1 0 48496 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_425
timestamp 1663859327
transform 1 0 48944 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_428
timestamp 1663859327
transform 1 0 49280 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_492
timestamp 1663859327
transform 1 0 56448 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_496
timestamp 1663859327
transform 1 0 56896 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_499
timestamp 1663859327
transform 1 0 57232 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_563
timestamp 1663859327
transform 1 0 64400 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_567
timestamp 1663859327
transform 1 0 64848 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_570
timestamp 1663859327
transform 1 0 65184 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_634
timestamp 1663859327
transform 1 0 72352 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_638
timestamp 1663859327
transform 1 0 72800 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_641
timestamp 1663859327
transform 1 0 73136 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_705
timestamp 1663859327
transform 1 0 80304 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_709
timestamp 1663859327
transform 1 0 80752 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_712
timestamp 1663859327
transform 1 0 81088 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_776
timestamp 1663859327
transform 1 0 88256 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_780
timestamp 1663859327
transform 1 0 88704 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_783
timestamp 1663859327
transform 1 0 89040 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_847
timestamp 1663859327
transform 1 0 96208 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_851
timestamp 1663859327
transform 1 0 96656 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_854
timestamp 1663859327
transform 1 0 96992 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_918
timestamp 1663859327
transform 1 0 104160 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_922
timestamp 1663859327
transform 1 0 104608 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_925
timestamp 1663859327
transform 1 0 104944 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_989
timestamp 1663859327
transform 1 0 112112 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_993
timestamp 1663859327
transform 1 0 112560 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_996
timestamp 1663859327
transform 1 0 112896 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_1028
timestamp 1663859327
transform 1 0 116480 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_1036
timestamp 1663859327
transform 1 0 117376 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_1044
timestamp 1663859327
transform 1 0 118272 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_2
timestamp 1663859327
transform 1 0 1568 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_7
timestamp 1663859327
transform 1 0 2128 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_23
timestamp 1663859327
transform 1 0 3920 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_31
timestamp 1663859327
transform 1 0 4816 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_37
timestamp 1663859327
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_101
timestamp 1663859327
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1663859327
transform 1 0 13104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_108
timestamp 1663859327
transform 1 0 13440 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_172
timestamp 1663859327
transform 1 0 20608 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_176
timestamp 1663859327
transform 1 0 21056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_179
timestamp 1663859327
transform 1 0 21392 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_243
timestamp 1663859327
transform 1 0 28560 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_247
timestamp 1663859327
transform 1 0 29008 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1663859327
transform 1 0 29344 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_314
timestamp 1663859327
transform 1 0 36512 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1663859327
transform 1 0 36960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1663859327
transform 1 0 37296 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_385
timestamp 1663859327
transform 1 0 44464 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1663859327
transform 1 0 44912 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_392
timestamp 1663859327
transform 1 0 45248 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_456
timestamp 1663859327
transform 1 0 52416 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_460
timestamp 1663859327
transform 1 0 52864 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_463
timestamp 1663859327
transform 1 0 53200 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_527
timestamp 1663859327
transform 1 0 60368 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_531
timestamp 1663859327
transform 1 0 60816 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_534
timestamp 1663859327
transform 1 0 61152 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_598
timestamp 1663859327
transform 1 0 68320 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_602
timestamp 1663859327
transform 1 0 68768 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_605
timestamp 1663859327
transform 1 0 69104 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_669
timestamp 1663859327
transform 1 0 76272 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_673
timestamp 1663859327
transform 1 0 76720 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_676
timestamp 1663859327
transform 1 0 77056 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_740
timestamp 1663859327
transform 1 0 84224 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_744
timestamp 1663859327
transform 1 0 84672 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_747
timestamp 1663859327
transform 1 0 85008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_811
timestamp 1663859327
transform 1 0 92176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_815
timestamp 1663859327
transform 1 0 92624 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_818
timestamp 1663859327
transform 1 0 92960 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_882
timestamp 1663859327
transform 1 0 100128 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_886
timestamp 1663859327
transform 1 0 100576 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_889
timestamp 1663859327
transform 1 0 100912 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_953
timestamp 1663859327
transform 1 0 108080 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_957
timestamp 1663859327
transform 1 0 108528 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_960
timestamp 1663859327
transform 1 0 108864 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1024
timestamp 1663859327
transform 1 0 116032 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_1028
timestamp 1663859327
transform 1 0 116480 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_1031
timestamp 1663859327
transform 1 0 116816 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_1039
timestamp 1663859327
transform 1 0 117712 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_1043
timestamp 1663859327
transform 1 0 118160 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_2
timestamp 1663859327
transform 1 0 1568 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_66
timestamp 1663859327
transform 1 0 8736 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_70
timestamp 1663859327
transform 1 0 9184 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_73
timestamp 1663859327
transform 1 0 9520 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_137
timestamp 1663859327
transform 1 0 16688 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_141
timestamp 1663859327
transform 1 0 17136 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_144
timestamp 1663859327
transform 1 0 17472 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_208
timestamp 1663859327
transform 1 0 24640 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1663859327
transform 1 0 25088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_215
timestamp 1663859327
transform 1 0 25424 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_279
timestamp 1663859327
transform 1 0 32592 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1663859327
transform 1 0 33040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1663859327
transform 1 0 33376 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_350
timestamp 1663859327
transform 1 0 40544 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1663859327
transform 1 0 40992 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_357
timestamp 1663859327
transform 1 0 41328 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_421
timestamp 1663859327
transform 1 0 48496 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_425
timestamp 1663859327
transform 1 0 48944 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_428
timestamp 1663859327
transform 1 0 49280 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_492
timestamp 1663859327
transform 1 0 56448 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_496
timestamp 1663859327
transform 1 0 56896 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_499
timestamp 1663859327
transform 1 0 57232 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_563
timestamp 1663859327
transform 1 0 64400 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_567
timestamp 1663859327
transform 1 0 64848 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_570
timestamp 1663859327
transform 1 0 65184 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_634
timestamp 1663859327
transform 1 0 72352 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_638
timestamp 1663859327
transform 1 0 72800 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_641
timestamp 1663859327
transform 1 0 73136 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_705
timestamp 1663859327
transform 1 0 80304 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_709
timestamp 1663859327
transform 1 0 80752 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_712
timestamp 1663859327
transform 1 0 81088 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_776
timestamp 1663859327
transform 1 0 88256 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_780
timestamp 1663859327
transform 1 0 88704 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_783
timestamp 1663859327
transform 1 0 89040 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_847
timestamp 1663859327
transform 1 0 96208 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_851
timestamp 1663859327
transform 1 0 96656 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_854
timestamp 1663859327
transform 1 0 96992 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_918
timestamp 1663859327
transform 1 0 104160 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_922
timestamp 1663859327
transform 1 0 104608 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_925
timestamp 1663859327
transform 1 0 104944 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_989
timestamp 1663859327
transform 1 0 112112 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_993
timestamp 1663859327
transform 1 0 112560 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_996
timestamp 1663859327
transform 1 0 112896 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_1028
timestamp 1663859327
transform 1 0 116480 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_1044
timestamp 1663859327
transform 1 0 118272 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_2
timestamp 1663859327
transform 1 0 1568 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_34
timestamp 1663859327
transform 1 0 5152 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_37
timestamp 1663859327
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_101
timestamp 1663859327
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1663859327
transform 1 0 13104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_108
timestamp 1663859327
transform 1 0 13440 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_172
timestamp 1663859327
transform 1 0 20608 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1663859327
transform 1 0 21056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_179
timestamp 1663859327
transform 1 0 21392 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_243
timestamp 1663859327
transform 1 0 28560 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1663859327
transform 1 0 29008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_250
timestamp 1663859327
transform 1 0 29344 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_314
timestamp 1663859327
transform 1 0 36512 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_318
timestamp 1663859327
transform 1 0 36960 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1663859327
transform 1 0 37296 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_385
timestamp 1663859327
transform 1 0 44464 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1663859327
transform 1 0 44912 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_392
timestamp 1663859327
transform 1 0 45248 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_456
timestamp 1663859327
transform 1 0 52416 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_460
timestamp 1663859327
transform 1 0 52864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_463
timestamp 1663859327
transform 1 0 53200 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_527
timestamp 1663859327
transform 1 0 60368 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_531
timestamp 1663859327
transform 1 0 60816 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_534
timestamp 1663859327
transform 1 0 61152 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_598
timestamp 1663859327
transform 1 0 68320 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_602
timestamp 1663859327
transform 1 0 68768 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_605
timestamp 1663859327
transform 1 0 69104 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_669
timestamp 1663859327
transform 1 0 76272 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_673
timestamp 1663859327
transform 1 0 76720 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_676
timestamp 1663859327
transform 1 0 77056 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_740
timestamp 1663859327
transform 1 0 84224 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_744
timestamp 1663859327
transform 1 0 84672 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_747
timestamp 1663859327
transform 1 0 85008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_811
timestamp 1663859327
transform 1 0 92176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_815
timestamp 1663859327
transform 1 0 92624 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_818
timestamp 1663859327
transform 1 0 92960 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_882
timestamp 1663859327
transform 1 0 100128 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_886
timestamp 1663859327
transform 1 0 100576 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_889
timestamp 1663859327
transform 1 0 100912 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_953
timestamp 1663859327
transform 1 0 108080 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_957
timestamp 1663859327
transform 1 0 108528 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_960
timestamp 1663859327
transform 1 0 108864 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1024
timestamp 1663859327
transform 1 0 116032 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_1028
timestamp 1663859327
transform 1 0 116480 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_1031
timestamp 1663859327
transform 1 0 116816 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_1039
timestamp 1663859327
transform 1 0 117712 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_1043
timestamp 1663859327
transform 1 0 118160 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_2
timestamp 1663859327
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_66
timestamp 1663859327
transform 1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_70
timestamp 1663859327
transform 1 0 9184 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_73
timestamp 1663859327
transform 1 0 9520 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_137
timestamp 1663859327
transform 1 0 16688 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1663859327
transform 1 0 17136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_144
timestamp 1663859327
transform 1 0 17472 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_208
timestamp 1663859327
transform 1 0 24640 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1663859327
transform 1 0 25088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_215
timestamp 1663859327
transform 1 0 25424 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_279
timestamp 1663859327
transform 1 0 32592 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_283
timestamp 1663859327
transform 1 0 33040 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1663859327
transform 1 0 33376 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_350
timestamp 1663859327
transform 1 0 40544 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1663859327
transform 1 0 40992 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_357
timestamp 1663859327
transform 1 0 41328 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_421
timestamp 1663859327
transform 1 0 48496 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_425
timestamp 1663859327
transform 1 0 48944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_428
timestamp 1663859327
transform 1 0 49280 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_492
timestamp 1663859327
transform 1 0 56448 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_496
timestamp 1663859327
transform 1 0 56896 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_499
timestamp 1663859327
transform 1 0 57232 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_563
timestamp 1663859327
transform 1 0 64400 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_567
timestamp 1663859327
transform 1 0 64848 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_570
timestamp 1663859327
transform 1 0 65184 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_634
timestamp 1663859327
transform 1 0 72352 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_638
timestamp 1663859327
transform 1 0 72800 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_641
timestamp 1663859327
transform 1 0 73136 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_705
timestamp 1663859327
transform 1 0 80304 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_709
timestamp 1663859327
transform 1 0 80752 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_712
timestamp 1663859327
transform 1 0 81088 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_776
timestamp 1663859327
transform 1 0 88256 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_780
timestamp 1663859327
transform 1 0 88704 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_783
timestamp 1663859327
transform 1 0 89040 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_847
timestamp 1663859327
transform 1 0 96208 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_851
timestamp 1663859327
transform 1 0 96656 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_854
timestamp 1663859327
transform 1 0 96992 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_918
timestamp 1663859327
transform 1 0 104160 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_922
timestamp 1663859327
transform 1 0 104608 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_925
timestamp 1663859327
transform 1 0 104944 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_989
timestamp 1663859327
transform 1 0 112112 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_993
timestamp 1663859327
transform 1 0 112560 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_996
timestamp 1663859327
transform 1 0 112896 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_1028
timestamp 1663859327
transform 1 0 116480 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_1044
timestamp 1663859327
transform 1 0 118272 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_2
timestamp 1663859327
transform 1 0 1568 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_7
timestamp 1663859327
transform 1 0 2128 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_23
timestamp 1663859327
transform 1 0 3920 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_31
timestamp 1663859327
transform 1 0 4816 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_37
timestamp 1663859327
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_101
timestamp 1663859327
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_105
timestamp 1663859327
transform 1 0 13104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_108
timestamp 1663859327
transform 1 0 13440 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_172
timestamp 1663859327
transform 1 0 20608 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_176
timestamp 1663859327
transform 1 0 21056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_179
timestamp 1663859327
transform 1 0 21392 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_243
timestamp 1663859327
transform 1 0 28560 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_247
timestamp 1663859327
transform 1 0 29008 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_250
timestamp 1663859327
transform 1 0 29344 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_314
timestamp 1663859327
transform 1 0 36512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1663859327
transform 1 0 36960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1663859327
transform 1 0 37296 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_385
timestamp 1663859327
transform 1 0 44464 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1663859327
transform 1 0 44912 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_392
timestamp 1663859327
transform 1 0 45248 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_456
timestamp 1663859327
transform 1 0 52416 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_460
timestamp 1663859327
transform 1 0 52864 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_463
timestamp 1663859327
transform 1 0 53200 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_527
timestamp 1663859327
transform 1 0 60368 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_531
timestamp 1663859327
transform 1 0 60816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_534
timestamp 1663859327
transform 1 0 61152 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_598
timestamp 1663859327
transform 1 0 68320 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_602
timestamp 1663859327
transform 1 0 68768 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_605
timestamp 1663859327
transform 1 0 69104 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_669
timestamp 1663859327
transform 1 0 76272 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_673
timestamp 1663859327
transform 1 0 76720 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_676
timestamp 1663859327
transform 1 0 77056 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_740
timestamp 1663859327
transform 1 0 84224 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_744
timestamp 1663859327
transform 1 0 84672 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_747
timestamp 1663859327
transform 1 0 85008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_811
timestamp 1663859327
transform 1 0 92176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_815
timestamp 1663859327
transform 1 0 92624 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_818
timestamp 1663859327
transform 1 0 92960 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_882
timestamp 1663859327
transform 1 0 100128 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_886
timestamp 1663859327
transform 1 0 100576 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_889
timestamp 1663859327
transform 1 0 100912 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_953
timestamp 1663859327
transform 1 0 108080 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_957
timestamp 1663859327
transform 1 0 108528 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_960
timestamp 1663859327
transform 1 0 108864 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1024
timestamp 1663859327
transform 1 0 116032 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_1028
timestamp 1663859327
transform 1 0 116480 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_1031
timestamp 1663859327
transform 1 0 116816 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_1039
timestamp 1663859327
transform 1 0 117712 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_1043
timestamp 1663859327
transform 1 0 118160 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_2
timestamp 1663859327
transform 1 0 1568 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_5
timestamp 1663859327
transform 1 0 1904 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_69
timestamp 1663859327
transform 1 0 9072 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_73
timestamp 1663859327
transform 1 0 9520 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_137
timestamp 1663859327
transform 1 0 16688 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_141
timestamp 1663859327
transform 1 0 17136 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_144
timestamp 1663859327
transform 1 0 17472 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_208
timestamp 1663859327
transform 1 0 24640 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1663859327
transform 1 0 25088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_215
timestamp 1663859327
transform 1 0 25424 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_279
timestamp 1663859327
transform 1 0 32592 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1663859327
transform 1 0 33040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1663859327
transform 1 0 33376 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_350
timestamp 1663859327
transform 1 0 40544 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1663859327
transform 1 0 40992 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_357
timestamp 1663859327
transform 1 0 41328 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_421
timestamp 1663859327
transform 1 0 48496 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_425
timestamp 1663859327
transform 1 0 48944 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_428
timestamp 1663859327
transform 1 0 49280 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_492
timestamp 1663859327
transform 1 0 56448 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_496
timestamp 1663859327
transform 1 0 56896 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_499
timestamp 1663859327
transform 1 0 57232 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_563
timestamp 1663859327
transform 1 0 64400 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_567
timestamp 1663859327
transform 1 0 64848 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_570
timestamp 1663859327
transform 1 0 65184 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_634
timestamp 1663859327
transform 1 0 72352 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_638
timestamp 1663859327
transform 1 0 72800 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_641
timestamp 1663859327
transform 1 0 73136 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_705
timestamp 1663859327
transform 1 0 80304 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_709
timestamp 1663859327
transform 1 0 80752 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_712
timestamp 1663859327
transform 1 0 81088 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_776
timestamp 1663859327
transform 1 0 88256 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_780
timestamp 1663859327
transform 1 0 88704 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_783
timestamp 1663859327
transform 1 0 89040 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_847
timestamp 1663859327
transform 1 0 96208 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_851
timestamp 1663859327
transform 1 0 96656 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_854
timestamp 1663859327
transform 1 0 96992 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_918
timestamp 1663859327
transform 1 0 104160 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_922
timestamp 1663859327
transform 1 0 104608 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_925
timestamp 1663859327
transform 1 0 104944 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_989
timestamp 1663859327
transform 1 0 112112 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_993
timestamp 1663859327
transform 1 0 112560 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_996
timestamp 1663859327
transform 1 0 112896 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_1028
timestamp 1663859327
transform 1 0 116480 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_1044
timestamp 1663859327
transform 1 0 118272 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_2
timestamp 1663859327
transform 1 0 1568 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_9
timestamp 1663859327
transform 1 0 2352 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_25
timestamp 1663859327
transform 1 0 4144 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_33
timestamp 1663859327
transform 1 0 5040 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_37
timestamp 1663859327
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_101
timestamp 1663859327
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_105
timestamp 1663859327
transform 1 0 13104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_108
timestamp 1663859327
transform 1 0 13440 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_172
timestamp 1663859327
transform 1 0 20608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_176
timestamp 1663859327
transform 1 0 21056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_179
timestamp 1663859327
transform 1 0 21392 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_243
timestamp 1663859327
transform 1 0 28560 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_247
timestamp 1663859327
transform 1 0 29008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_250
timestamp 1663859327
transform 1 0 29344 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_314
timestamp 1663859327
transform 1 0 36512 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_318
timestamp 1663859327
transform 1 0 36960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_321
timestamp 1663859327
transform 1 0 37296 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_385
timestamp 1663859327
transform 1 0 44464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_389
timestamp 1663859327
transform 1 0 44912 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_392
timestamp 1663859327
transform 1 0 45248 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_456
timestamp 1663859327
transform 1 0 52416 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_460
timestamp 1663859327
transform 1 0 52864 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_463
timestamp 1663859327
transform 1 0 53200 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_527
timestamp 1663859327
transform 1 0 60368 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_531
timestamp 1663859327
transform 1 0 60816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_534
timestamp 1663859327
transform 1 0 61152 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_598
timestamp 1663859327
transform 1 0 68320 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_602
timestamp 1663859327
transform 1 0 68768 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_605
timestamp 1663859327
transform 1 0 69104 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_669
timestamp 1663859327
transform 1 0 76272 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_673
timestamp 1663859327
transform 1 0 76720 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_676
timestamp 1663859327
transform 1 0 77056 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_740
timestamp 1663859327
transform 1 0 84224 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_744
timestamp 1663859327
transform 1 0 84672 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_747
timestamp 1663859327
transform 1 0 85008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_811
timestamp 1663859327
transform 1 0 92176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_815
timestamp 1663859327
transform 1 0 92624 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_818
timestamp 1663859327
transform 1 0 92960 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_882
timestamp 1663859327
transform 1 0 100128 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_886
timestamp 1663859327
transform 1 0 100576 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_889
timestamp 1663859327
transform 1 0 100912 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_953
timestamp 1663859327
transform 1 0 108080 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_957
timestamp 1663859327
transform 1 0 108528 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_960
timestamp 1663859327
transform 1 0 108864 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1024
timestamp 1663859327
transform 1 0 116032 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_1028
timestamp 1663859327
transform 1 0 116480 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_1031
timestamp 1663859327
transform 1 0 116816 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_1039
timestamp 1663859327
transform 1 0 117712 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_1043
timestamp 1663859327
transform 1 0 118160 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_2
timestamp 1663859327
transform 1 0 1568 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_42
timestamp 1663859327
transform 1 0 6048 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_46
timestamp 1663859327
transform 1 0 6496 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_62
timestamp 1663859327
transform 1 0 8288 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_70
timestamp 1663859327
transform 1 0 9184 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_73
timestamp 1663859327
transform 1 0 9520 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_137
timestamp 1663859327
transform 1 0 16688 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_141
timestamp 1663859327
transform 1 0 17136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_144
timestamp 1663859327
transform 1 0 17472 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_208
timestamp 1663859327
transform 1 0 24640 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_212
timestamp 1663859327
transform 1 0 25088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_215
timestamp 1663859327
transform 1 0 25424 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_279
timestamp 1663859327
transform 1 0 32592 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_283
timestamp 1663859327
transform 1 0 33040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_286
timestamp 1663859327
transform 1 0 33376 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_350
timestamp 1663859327
transform 1 0 40544 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_354
timestamp 1663859327
transform 1 0 40992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_357
timestamp 1663859327
transform 1 0 41328 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_421
timestamp 1663859327
transform 1 0 48496 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_425
timestamp 1663859327
transform 1 0 48944 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_428
timestamp 1663859327
transform 1 0 49280 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_492
timestamp 1663859327
transform 1 0 56448 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_496
timestamp 1663859327
transform 1 0 56896 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_499
timestamp 1663859327
transform 1 0 57232 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_563
timestamp 1663859327
transform 1 0 64400 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_567
timestamp 1663859327
transform 1 0 64848 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_570
timestamp 1663859327
transform 1 0 65184 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_634
timestamp 1663859327
transform 1 0 72352 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_638
timestamp 1663859327
transform 1 0 72800 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_641
timestamp 1663859327
transform 1 0 73136 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_705
timestamp 1663859327
transform 1 0 80304 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_709
timestamp 1663859327
transform 1 0 80752 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_712
timestamp 1663859327
transform 1 0 81088 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_776
timestamp 1663859327
transform 1 0 88256 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_780
timestamp 1663859327
transform 1 0 88704 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_783
timestamp 1663859327
transform 1 0 89040 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_847
timestamp 1663859327
transform 1 0 96208 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_851
timestamp 1663859327
transform 1 0 96656 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_854
timestamp 1663859327
transform 1 0 96992 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_918
timestamp 1663859327
transform 1 0 104160 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_922
timestamp 1663859327
transform 1 0 104608 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_925
timestamp 1663859327
transform 1 0 104944 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_989
timestamp 1663859327
transform 1 0 112112 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_993
timestamp 1663859327
transform 1 0 112560 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_996
timestamp 1663859327
transform 1 0 112896 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_1028
timestamp 1663859327
transform 1 0 116480 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_1044
timestamp 1663859327
transform 1 0 118272 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_2
timestamp 1663859327
transform 1 0 1568 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_4
timestamp 1663859327
transform 1 0 1792 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_7
timestamp 1663859327
transform 1 0 2128 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_15
timestamp 1663859327
transform 1 0 3024 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_22
timestamp 1663859327
transform 1 0 3808 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_26
timestamp 1663859327
transform 1 0 4256 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_34
timestamp 1663859327
transform 1 0 5152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_37
timestamp 1663859327
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_101
timestamp 1663859327
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_105
timestamp 1663859327
transform 1 0 13104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_108
timestamp 1663859327
transform 1 0 13440 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_172
timestamp 1663859327
transform 1 0 20608 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_176
timestamp 1663859327
transform 1 0 21056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_179
timestamp 1663859327
transform 1 0 21392 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_243
timestamp 1663859327
transform 1 0 28560 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_247
timestamp 1663859327
transform 1 0 29008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_250
timestamp 1663859327
transform 1 0 29344 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_314
timestamp 1663859327
transform 1 0 36512 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_318
timestamp 1663859327
transform 1 0 36960 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_321
timestamp 1663859327
transform 1 0 37296 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_385
timestamp 1663859327
transform 1 0 44464 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_389
timestamp 1663859327
transform 1 0 44912 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_392
timestamp 1663859327
transform 1 0 45248 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_456
timestamp 1663859327
transform 1 0 52416 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_460
timestamp 1663859327
transform 1 0 52864 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_463
timestamp 1663859327
transform 1 0 53200 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_495
timestamp 1663859327
transform 1 0 56784 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_511
timestamp 1663859327
transform 1 0 58576 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_515
timestamp 1663859327
transform 1 0 59024 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_522
timestamp 1663859327
transform 1 0 59808 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_526
timestamp 1663859327
transform 1 0 60256 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_530
timestamp 1663859327
transform 1 0 60704 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_534
timestamp 1663859327
transform 1 0 61152 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_598
timestamp 1663859327
transform 1 0 68320 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_602
timestamp 1663859327
transform 1 0 68768 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_605
timestamp 1663859327
transform 1 0 69104 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_669
timestamp 1663859327
transform 1 0 76272 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_673
timestamp 1663859327
transform 1 0 76720 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_676
timestamp 1663859327
transform 1 0 77056 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_740
timestamp 1663859327
transform 1 0 84224 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_744
timestamp 1663859327
transform 1 0 84672 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_747
timestamp 1663859327
transform 1 0 85008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_811
timestamp 1663859327
transform 1 0 92176 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_815
timestamp 1663859327
transform 1 0 92624 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_818
timestamp 1663859327
transform 1 0 92960 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_882
timestamp 1663859327
transform 1 0 100128 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_886
timestamp 1663859327
transform 1 0 100576 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_889
timestamp 1663859327
transform 1 0 100912 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_953
timestamp 1663859327
transform 1 0 108080 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_957
timestamp 1663859327
transform 1 0 108528 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_960
timestamp 1663859327
transform 1 0 108864 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_1024
timestamp 1663859327
transform 1 0 116032 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1028
timestamp 1663859327
transform 1 0 116480 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_1031
timestamp 1663859327
transform 1 0 116816 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1039
timestamp 1663859327
transform 1 0 117712 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_1044
timestamp 1663859327
transform 1 0 118272 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_2
timestamp 1663859327
transform 1 0 1568 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_14
timestamp 1663859327
transform 1 0 2912 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_18
timestamp 1663859327
transform 1 0 3360 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_50
timestamp 1663859327
transform 1 0 6944 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_66
timestamp 1663859327
transform 1 0 8736 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_70
timestamp 1663859327
transform 1 0 9184 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_73
timestamp 1663859327
transform 1 0 9520 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_137
timestamp 1663859327
transform 1 0 16688 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_141
timestamp 1663859327
transform 1 0 17136 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_144
timestamp 1663859327
transform 1 0 17472 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_160
timestamp 1663859327
transform 1 0 19264 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_164
timestamp 1663859327
transform 1 0 19712 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_169
timestamp 1663859327
transform 1 0 20272 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_173
timestamp 1663859327
transform 1 0 20720 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_205
timestamp 1663859327
transform 1 0 24304 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_215
timestamp 1663859327
transform 1 0 25424 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_279
timestamp 1663859327
transform 1 0 32592 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_283
timestamp 1663859327
transform 1 0 33040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_286
timestamp 1663859327
transform 1 0 33376 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_350
timestamp 1663859327
transform 1 0 40544 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_354
timestamp 1663859327
transform 1 0 40992 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_357
timestamp 1663859327
transform 1 0 41328 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_421
timestamp 1663859327
transform 1 0 48496 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_425
timestamp 1663859327
transform 1 0 48944 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_428
timestamp 1663859327
transform 1 0 49280 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_492
timestamp 1663859327
transform 1 0 56448 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_496
timestamp 1663859327
transform 1 0 56896 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_499
timestamp 1663859327
transform 1 0 57232 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_563
timestamp 1663859327
transform 1 0 64400 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_567
timestamp 1663859327
transform 1 0 64848 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_570
timestamp 1663859327
transform 1 0 65184 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_634
timestamp 1663859327
transform 1 0 72352 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_638
timestamp 1663859327
transform 1 0 72800 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_641
timestamp 1663859327
transform 1 0 73136 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_705
timestamp 1663859327
transform 1 0 80304 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_709
timestamp 1663859327
transform 1 0 80752 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_712
timestamp 1663859327
transform 1 0 81088 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_776
timestamp 1663859327
transform 1 0 88256 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_780
timestamp 1663859327
transform 1 0 88704 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_783
timestamp 1663859327
transform 1 0 89040 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_847
timestamp 1663859327
transform 1 0 96208 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_851
timestamp 1663859327
transform 1 0 96656 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_854
timestamp 1663859327
transform 1 0 96992 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_918
timestamp 1663859327
transform 1 0 104160 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_922
timestamp 1663859327
transform 1 0 104608 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_925
timestamp 1663859327
transform 1 0 104944 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_989
timestamp 1663859327
transform 1 0 112112 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_993
timestamp 1663859327
transform 1 0 112560 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_996
timestamp 1663859327
transform 1 0 112896 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_1028
timestamp 1663859327
transform 1 0 116480 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_1036
timestamp 1663859327
transform 1 0 117376 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_1044
timestamp 1663859327
transform 1 0 118272 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_2
timestamp 1663859327
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_34
timestamp 1663859327
transform 1 0 5152 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_37
timestamp 1663859327
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_101
timestamp 1663859327
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_105
timestamp 1663859327
transform 1 0 13104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_108
timestamp 1663859327
transform 1 0 13440 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_172
timestamp 1663859327
transform 1 0 20608 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_176
timestamp 1663859327
transform 1 0 21056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_179
timestamp 1663859327
transform 1 0 21392 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_243
timestamp 1663859327
transform 1 0 28560 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_247
timestamp 1663859327
transform 1 0 29008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_250
timestamp 1663859327
transform 1 0 29344 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_314
timestamp 1663859327
transform 1 0 36512 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_318
timestamp 1663859327
transform 1 0 36960 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_321
timestamp 1663859327
transform 1 0 37296 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_385
timestamp 1663859327
transform 1 0 44464 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_389
timestamp 1663859327
transform 1 0 44912 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_392
timestamp 1663859327
transform 1 0 45248 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_456
timestamp 1663859327
transform 1 0 52416 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_460
timestamp 1663859327
transform 1 0 52864 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_463
timestamp 1663859327
transform 1 0 53200 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_527
timestamp 1663859327
transform 1 0 60368 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_531
timestamp 1663859327
transform 1 0 60816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_534
timestamp 1663859327
transform 1 0 61152 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_598
timestamp 1663859327
transform 1 0 68320 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_602
timestamp 1663859327
transform 1 0 68768 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_605
timestamp 1663859327
transform 1 0 69104 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_669
timestamp 1663859327
transform 1 0 76272 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_673
timestamp 1663859327
transform 1 0 76720 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_676
timestamp 1663859327
transform 1 0 77056 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_740
timestamp 1663859327
transform 1 0 84224 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_744
timestamp 1663859327
transform 1 0 84672 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_747
timestamp 1663859327
transform 1 0 85008 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_811
timestamp 1663859327
transform 1 0 92176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_815
timestamp 1663859327
transform 1 0 92624 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_818
timestamp 1663859327
transform 1 0 92960 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_882
timestamp 1663859327
transform 1 0 100128 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_886
timestamp 1663859327
transform 1 0 100576 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_889
timestamp 1663859327
transform 1 0 100912 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_953
timestamp 1663859327
transform 1 0 108080 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_957
timestamp 1663859327
transform 1 0 108528 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_960
timestamp 1663859327
transform 1 0 108864 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_1024
timestamp 1663859327
transform 1 0 116032 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1028
timestamp 1663859327
transform 1 0 116480 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_1031
timestamp 1663859327
transform 1 0 116816 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1039
timestamp 1663859327
transform 1 0 117712 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_1044
timestamp 1663859327
transform 1 0 118272 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_2
timestamp 1663859327
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_66
timestamp 1663859327
transform 1 0 8736 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_70
timestamp 1663859327
transform 1 0 9184 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_73
timestamp 1663859327
transform 1 0 9520 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_137
timestamp 1663859327
transform 1 0 16688 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_141
timestamp 1663859327
transform 1 0 17136 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_144
timestamp 1663859327
transform 1 0 17472 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_208
timestamp 1663859327
transform 1 0 24640 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_212
timestamp 1663859327
transform 1 0 25088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_215
timestamp 1663859327
transform 1 0 25424 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_279
timestamp 1663859327
transform 1 0 32592 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_283
timestamp 1663859327
transform 1 0 33040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_286
timestamp 1663859327
transform 1 0 33376 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_350
timestamp 1663859327
transform 1 0 40544 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_354
timestamp 1663859327
transform 1 0 40992 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_357
timestamp 1663859327
transform 1 0 41328 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_421
timestamp 1663859327
transform 1 0 48496 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_425
timestamp 1663859327
transform 1 0 48944 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_428
timestamp 1663859327
transform 1 0 49280 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_492
timestamp 1663859327
transform 1 0 56448 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_496
timestamp 1663859327
transform 1 0 56896 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_499
timestamp 1663859327
transform 1 0 57232 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_563
timestamp 1663859327
transform 1 0 64400 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_567
timestamp 1663859327
transform 1 0 64848 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_570
timestamp 1663859327
transform 1 0 65184 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_634
timestamp 1663859327
transform 1 0 72352 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_638
timestamp 1663859327
transform 1 0 72800 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_641
timestamp 1663859327
transform 1 0 73136 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_705
timestamp 1663859327
transform 1 0 80304 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_709
timestamp 1663859327
transform 1 0 80752 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_712
timestamp 1663859327
transform 1 0 81088 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_776
timestamp 1663859327
transform 1 0 88256 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_780
timestamp 1663859327
transform 1 0 88704 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_783
timestamp 1663859327
transform 1 0 89040 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_847
timestamp 1663859327
transform 1 0 96208 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_851
timestamp 1663859327
transform 1 0 96656 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_854
timestamp 1663859327
transform 1 0 96992 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_918
timestamp 1663859327
transform 1 0 104160 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_922
timestamp 1663859327
transform 1 0 104608 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_925
timestamp 1663859327
transform 1 0 104944 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_989
timestamp 1663859327
transform 1 0 112112 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_993
timestamp 1663859327
transform 1 0 112560 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_996
timestamp 1663859327
transform 1 0 112896 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_1028
timestamp 1663859327
transform 1 0 116480 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_1044
timestamp 1663859327
transform 1 0 118272 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_86_2
timestamp 1663859327
transform 1 0 1568 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_34
timestamp 1663859327
transform 1 0 5152 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_37
timestamp 1663859327
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_101
timestamp 1663859327
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_105
timestamp 1663859327
transform 1 0 13104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_108
timestamp 1663859327
transform 1 0 13440 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_172
timestamp 1663859327
transform 1 0 20608 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_176
timestamp 1663859327
transform 1 0 21056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_179
timestamp 1663859327
transform 1 0 21392 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_243
timestamp 1663859327
transform 1 0 28560 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_247
timestamp 1663859327
transform 1 0 29008 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_250
timestamp 1663859327
transform 1 0 29344 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_314
timestamp 1663859327
transform 1 0 36512 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_318
timestamp 1663859327
transform 1 0 36960 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_321
timestamp 1663859327
transform 1 0 37296 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_385
timestamp 1663859327
transform 1 0 44464 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_389
timestamp 1663859327
transform 1 0 44912 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_392
timestamp 1663859327
transform 1 0 45248 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_456
timestamp 1663859327
transform 1 0 52416 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_460
timestamp 1663859327
transform 1 0 52864 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_463
timestamp 1663859327
transform 1 0 53200 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_527
timestamp 1663859327
transform 1 0 60368 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_531
timestamp 1663859327
transform 1 0 60816 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_534
timestamp 1663859327
transform 1 0 61152 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_598
timestamp 1663859327
transform 1 0 68320 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_602
timestamp 1663859327
transform 1 0 68768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_605
timestamp 1663859327
transform 1 0 69104 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_669
timestamp 1663859327
transform 1 0 76272 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_673
timestamp 1663859327
transform 1 0 76720 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_676
timestamp 1663859327
transform 1 0 77056 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_740
timestamp 1663859327
transform 1 0 84224 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_744
timestamp 1663859327
transform 1 0 84672 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_747
timestamp 1663859327
transform 1 0 85008 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_811
timestamp 1663859327
transform 1 0 92176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_815
timestamp 1663859327
transform 1 0 92624 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_818
timestamp 1663859327
transform 1 0 92960 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_882
timestamp 1663859327
transform 1 0 100128 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_886
timestamp 1663859327
transform 1 0 100576 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_889
timestamp 1663859327
transform 1 0 100912 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_953
timestamp 1663859327
transform 1 0 108080 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_957
timestamp 1663859327
transform 1 0 108528 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_960
timestamp 1663859327
transform 1 0 108864 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1024
timestamp 1663859327
transform 1 0 116032 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_1028
timestamp 1663859327
transform 1 0 116480 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_1031
timestamp 1663859327
transform 1 0 116816 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_1039
timestamp 1663859327
transform 1 0 117712 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_1043
timestamp 1663859327
transform 1 0 118160 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_2
timestamp 1663859327
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_66
timestamp 1663859327
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_70
timestamp 1663859327
transform 1 0 9184 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_73
timestamp 1663859327
transform 1 0 9520 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_137
timestamp 1663859327
transform 1 0 16688 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_141
timestamp 1663859327
transform 1 0 17136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_144
timestamp 1663859327
transform 1 0 17472 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_208
timestamp 1663859327
transform 1 0 24640 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_212
timestamp 1663859327
transform 1 0 25088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_215
timestamp 1663859327
transform 1 0 25424 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_279
timestamp 1663859327
transform 1 0 32592 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_283
timestamp 1663859327
transform 1 0 33040 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_286
timestamp 1663859327
transform 1 0 33376 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_350
timestamp 1663859327
transform 1 0 40544 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_354
timestamp 1663859327
transform 1 0 40992 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_357
timestamp 1663859327
transform 1 0 41328 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_421
timestamp 1663859327
transform 1 0 48496 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_425
timestamp 1663859327
transform 1 0 48944 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_428
timestamp 1663859327
transform 1 0 49280 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_492
timestamp 1663859327
transform 1 0 56448 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_496
timestamp 1663859327
transform 1 0 56896 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_499
timestamp 1663859327
transform 1 0 57232 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_563
timestamp 1663859327
transform 1 0 64400 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_567
timestamp 1663859327
transform 1 0 64848 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_570
timestamp 1663859327
transform 1 0 65184 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_634
timestamp 1663859327
transform 1 0 72352 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_638
timestamp 1663859327
transform 1 0 72800 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_641
timestamp 1663859327
transform 1 0 73136 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_705
timestamp 1663859327
transform 1 0 80304 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_709
timestamp 1663859327
transform 1 0 80752 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_712
timestamp 1663859327
transform 1 0 81088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_776
timestamp 1663859327
transform 1 0 88256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_780
timestamp 1663859327
transform 1 0 88704 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_783
timestamp 1663859327
transform 1 0 89040 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_847
timestamp 1663859327
transform 1 0 96208 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_851
timestamp 1663859327
transform 1 0 96656 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_854
timestamp 1663859327
transform 1 0 96992 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_918
timestamp 1663859327
transform 1 0 104160 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_922
timestamp 1663859327
transform 1 0 104608 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_925
timestamp 1663859327
transform 1 0 104944 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_989
timestamp 1663859327
transform 1 0 112112 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_993
timestamp 1663859327
transform 1 0 112560 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_996
timestamp 1663859327
transform 1 0 112896 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_1028
timestamp 1663859327
transform 1 0 116480 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_1044
timestamp 1663859327
transform 1 0 118272 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_2
timestamp 1663859327
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_34
timestamp 1663859327
transform 1 0 5152 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_37
timestamp 1663859327
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_101
timestamp 1663859327
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_105
timestamp 1663859327
transform 1 0 13104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_108
timestamp 1663859327
transform 1 0 13440 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_172
timestamp 1663859327
transform 1 0 20608 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_176
timestamp 1663859327
transform 1 0 21056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_179
timestamp 1663859327
transform 1 0 21392 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_243
timestamp 1663859327
transform 1 0 28560 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_247
timestamp 1663859327
transform 1 0 29008 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_250
timestamp 1663859327
transform 1 0 29344 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_314
timestamp 1663859327
transform 1 0 36512 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_318
timestamp 1663859327
transform 1 0 36960 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_321
timestamp 1663859327
transform 1 0 37296 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_385
timestamp 1663859327
transform 1 0 44464 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_389
timestamp 1663859327
transform 1 0 44912 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_392
timestamp 1663859327
transform 1 0 45248 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_456
timestamp 1663859327
transform 1 0 52416 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_460
timestamp 1663859327
transform 1 0 52864 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_463
timestamp 1663859327
transform 1 0 53200 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_527
timestamp 1663859327
transform 1 0 60368 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_531
timestamp 1663859327
transform 1 0 60816 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_534
timestamp 1663859327
transform 1 0 61152 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_598
timestamp 1663859327
transform 1 0 68320 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_602
timestamp 1663859327
transform 1 0 68768 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_605
timestamp 1663859327
transform 1 0 69104 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_669
timestamp 1663859327
transform 1 0 76272 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_673
timestamp 1663859327
transform 1 0 76720 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_676
timestamp 1663859327
transform 1 0 77056 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_740
timestamp 1663859327
transform 1 0 84224 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_744
timestamp 1663859327
transform 1 0 84672 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_747
timestamp 1663859327
transform 1 0 85008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_811
timestamp 1663859327
transform 1 0 92176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_815
timestamp 1663859327
transform 1 0 92624 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_818
timestamp 1663859327
transform 1 0 92960 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_882
timestamp 1663859327
transform 1 0 100128 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_886
timestamp 1663859327
transform 1 0 100576 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_889
timestamp 1663859327
transform 1 0 100912 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_953
timestamp 1663859327
transform 1 0 108080 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_957
timestamp 1663859327
transform 1 0 108528 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_960
timestamp 1663859327
transform 1 0 108864 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1024
timestamp 1663859327
transform 1 0 116032 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_1028
timestamp 1663859327
transform 1 0 116480 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_1031
timestamp 1663859327
transform 1 0 116816 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_1039
timestamp 1663859327
transform 1 0 117712 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_1043
timestamp 1663859327
transform 1 0 118160 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_2
timestamp 1663859327
transform 1 0 1568 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_7
timestamp 1663859327
transform 1 0 2128 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_73
timestamp 1663859327
transform 1 0 9520 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_137
timestamp 1663859327
transform 1 0 16688 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_141
timestamp 1663859327
transform 1 0 17136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_144
timestamp 1663859327
transform 1 0 17472 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_208
timestamp 1663859327
transform 1 0 24640 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_212
timestamp 1663859327
transform 1 0 25088 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_215
timestamp 1663859327
transform 1 0 25424 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_279
timestamp 1663859327
transform 1 0 32592 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_283
timestamp 1663859327
transform 1 0 33040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_286
timestamp 1663859327
transform 1 0 33376 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_350
timestamp 1663859327
transform 1 0 40544 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_354
timestamp 1663859327
transform 1 0 40992 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_357
timestamp 1663859327
transform 1 0 41328 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_421
timestamp 1663859327
transform 1 0 48496 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_425
timestamp 1663859327
transform 1 0 48944 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_428
timestamp 1663859327
transform 1 0 49280 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_492
timestamp 1663859327
transform 1 0 56448 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_496
timestamp 1663859327
transform 1 0 56896 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_499
timestamp 1663859327
transform 1 0 57232 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_563
timestamp 1663859327
transform 1 0 64400 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_567
timestamp 1663859327
transform 1 0 64848 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_570
timestamp 1663859327
transform 1 0 65184 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_634
timestamp 1663859327
transform 1 0 72352 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_638
timestamp 1663859327
transform 1 0 72800 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_641
timestamp 1663859327
transform 1 0 73136 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_705
timestamp 1663859327
transform 1 0 80304 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_709
timestamp 1663859327
transform 1 0 80752 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_712
timestamp 1663859327
transform 1 0 81088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_776
timestamp 1663859327
transform 1 0 88256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_780
timestamp 1663859327
transform 1 0 88704 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_783
timestamp 1663859327
transform 1 0 89040 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_847
timestamp 1663859327
transform 1 0 96208 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_851
timestamp 1663859327
transform 1 0 96656 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_854
timestamp 1663859327
transform 1 0 96992 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_918
timestamp 1663859327
transform 1 0 104160 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_922
timestamp 1663859327
transform 1 0 104608 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_925
timestamp 1663859327
transform 1 0 104944 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_989
timestamp 1663859327
transform 1 0 112112 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_993
timestamp 1663859327
transform 1 0 112560 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_996
timestamp 1663859327
transform 1 0 112896 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_1028
timestamp 1663859327
transform 1 0 116480 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_1044
timestamp 1663859327
transform 1 0 118272 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_2
timestamp 1663859327
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_34
timestamp 1663859327
transform 1 0 5152 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_37
timestamp 1663859327
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_101
timestamp 1663859327
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_105
timestamp 1663859327
transform 1 0 13104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_108
timestamp 1663859327
transform 1 0 13440 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_172
timestamp 1663859327
transform 1 0 20608 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_176
timestamp 1663859327
transform 1 0 21056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_179
timestamp 1663859327
transform 1 0 21392 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_243
timestamp 1663859327
transform 1 0 28560 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_247
timestamp 1663859327
transform 1 0 29008 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_250
timestamp 1663859327
transform 1 0 29344 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_314
timestamp 1663859327
transform 1 0 36512 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_318
timestamp 1663859327
transform 1 0 36960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_321
timestamp 1663859327
transform 1 0 37296 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_385
timestamp 1663859327
transform 1 0 44464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_389
timestamp 1663859327
transform 1 0 44912 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_392
timestamp 1663859327
transform 1 0 45248 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_456
timestamp 1663859327
transform 1 0 52416 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_460
timestamp 1663859327
transform 1 0 52864 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_463
timestamp 1663859327
transform 1 0 53200 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_527
timestamp 1663859327
transform 1 0 60368 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_531
timestamp 1663859327
transform 1 0 60816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_534
timestamp 1663859327
transform 1 0 61152 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_598
timestamp 1663859327
transform 1 0 68320 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_602
timestamp 1663859327
transform 1 0 68768 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_605
timestamp 1663859327
transform 1 0 69104 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_669
timestamp 1663859327
transform 1 0 76272 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_673
timestamp 1663859327
transform 1 0 76720 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_676
timestamp 1663859327
transform 1 0 77056 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_740
timestamp 1663859327
transform 1 0 84224 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_744
timestamp 1663859327
transform 1 0 84672 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_747
timestamp 1663859327
transform 1 0 85008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_811
timestamp 1663859327
transform 1 0 92176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_815
timestamp 1663859327
transform 1 0 92624 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_818
timestamp 1663859327
transform 1 0 92960 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_882
timestamp 1663859327
transform 1 0 100128 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_886
timestamp 1663859327
transform 1 0 100576 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_889
timestamp 1663859327
transform 1 0 100912 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_953
timestamp 1663859327
transform 1 0 108080 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_957
timestamp 1663859327
transform 1 0 108528 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_960
timestamp 1663859327
transform 1 0 108864 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_1024
timestamp 1663859327
transform 1 0 116032 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1028
timestamp 1663859327
transform 1 0 116480 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_1031
timestamp 1663859327
transform 1 0 116816 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1039
timestamp 1663859327
transform 1 0 117712 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_1044
timestamp 1663859327
transform 1 0 118272 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_2
timestamp 1663859327
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_66
timestamp 1663859327
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_70
timestamp 1663859327
transform 1 0 9184 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_73
timestamp 1663859327
transform 1 0 9520 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_137
timestamp 1663859327
transform 1 0 16688 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_141
timestamp 1663859327
transform 1 0 17136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_144
timestamp 1663859327
transform 1 0 17472 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_208
timestamp 1663859327
transform 1 0 24640 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_212
timestamp 1663859327
transform 1 0 25088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_215
timestamp 1663859327
transform 1 0 25424 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_279
timestamp 1663859327
transform 1 0 32592 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_283
timestamp 1663859327
transform 1 0 33040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_286
timestamp 1663859327
transform 1 0 33376 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_350
timestamp 1663859327
transform 1 0 40544 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_354
timestamp 1663859327
transform 1 0 40992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_357
timestamp 1663859327
transform 1 0 41328 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_421
timestamp 1663859327
transform 1 0 48496 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_425
timestamp 1663859327
transform 1 0 48944 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_428
timestamp 1663859327
transform 1 0 49280 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_492
timestamp 1663859327
transform 1 0 56448 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_496
timestamp 1663859327
transform 1 0 56896 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_499
timestamp 1663859327
transform 1 0 57232 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_563
timestamp 1663859327
transform 1 0 64400 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_567
timestamp 1663859327
transform 1 0 64848 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_570
timestamp 1663859327
transform 1 0 65184 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_634
timestamp 1663859327
transform 1 0 72352 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_638
timestamp 1663859327
transform 1 0 72800 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_641
timestamp 1663859327
transform 1 0 73136 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_705
timestamp 1663859327
transform 1 0 80304 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_709
timestamp 1663859327
transform 1 0 80752 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_712
timestamp 1663859327
transform 1 0 81088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_776
timestamp 1663859327
transform 1 0 88256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_780
timestamp 1663859327
transform 1 0 88704 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_783
timestamp 1663859327
transform 1 0 89040 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_847
timestamp 1663859327
transform 1 0 96208 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_851
timestamp 1663859327
transform 1 0 96656 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_854
timestamp 1663859327
transform 1 0 96992 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_918
timestamp 1663859327
transform 1 0 104160 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_922
timestamp 1663859327
transform 1 0 104608 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_925
timestamp 1663859327
transform 1 0 104944 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_989
timestamp 1663859327
transform 1 0 112112 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_993
timestamp 1663859327
transform 1 0 112560 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_996
timestamp 1663859327
transform 1 0 112896 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_1028
timestamp 1663859327
transform 1 0 116480 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_1044
timestamp 1663859327
transform 1 0 118272 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_2
timestamp 1663859327
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_34
timestamp 1663859327
transform 1 0 5152 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_37
timestamp 1663859327
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_101
timestamp 1663859327
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_105
timestamp 1663859327
transform 1 0 13104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_108
timestamp 1663859327
transform 1 0 13440 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_172
timestamp 1663859327
transform 1 0 20608 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_176
timestamp 1663859327
transform 1 0 21056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_179
timestamp 1663859327
transform 1 0 21392 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_243
timestamp 1663859327
transform 1 0 28560 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_247
timestamp 1663859327
transform 1 0 29008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_250
timestamp 1663859327
transform 1 0 29344 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_314
timestamp 1663859327
transform 1 0 36512 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_318
timestamp 1663859327
transform 1 0 36960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_321
timestamp 1663859327
transform 1 0 37296 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_385
timestamp 1663859327
transform 1 0 44464 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_389
timestamp 1663859327
transform 1 0 44912 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_392
timestamp 1663859327
transform 1 0 45248 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_456
timestamp 1663859327
transform 1 0 52416 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_460
timestamp 1663859327
transform 1 0 52864 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_463
timestamp 1663859327
transform 1 0 53200 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_527
timestamp 1663859327
transform 1 0 60368 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_531
timestamp 1663859327
transform 1 0 60816 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_534
timestamp 1663859327
transform 1 0 61152 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_598
timestamp 1663859327
transform 1 0 68320 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_602
timestamp 1663859327
transform 1 0 68768 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_605
timestamp 1663859327
transform 1 0 69104 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_669
timestamp 1663859327
transform 1 0 76272 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_673
timestamp 1663859327
transform 1 0 76720 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_676
timestamp 1663859327
transform 1 0 77056 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_740
timestamp 1663859327
transform 1 0 84224 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_744
timestamp 1663859327
transform 1 0 84672 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_747
timestamp 1663859327
transform 1 0 85008 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_811
timestamp 1663859327
transform 1 0 92176 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_815
timestamp 1663859327
transform 1 0 92624 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_818
timestamp 1663859327
transform 1 0 92960 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_882
timestamp 1663859327
transform 1 0 100128 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_886
timestamp 1663859327
transform 1 0 100576 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_889
timestamp 1663859327
transform 1 0 100912 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_953
timestamp 1663859327
transform 1 0 108080 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_957
timestamp 1663859327
transform 1 0 108528 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_960
timestamp 1663859327
transform 1 0 108864 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1024
timestamp 1663859327
transform 1 0 116032 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_1028
timestamp 1663859327
transform 1 0 116480 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_1031
timestamp 1663859327
transform 1 0 116816 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_1039
timestamp 1663859327
transform 1 0 117712 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_1043
timestamp 1663859327
transform 1 0 118160 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_2
timestamp 1663859327
transform 1 0 1568 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_66
timestamp 1663859327
transform 1 0 8736 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_70
timestamp 1663859327
transform 1 0 9184 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_73
timestamp 1663859327
transform 1 0 9520 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_137
timestamp 1663859327
transform 1 0 16688 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_141
timestamp 1663859327
transform 1 0 17136 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_144
timestamp 1663859327
transform 1 0 17472 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_208
timestamp 1663859327
transform 1 0 24640 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_212
timestamp 1663859327
transform 1 0 25088 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_215
timestamp 1663859327
transform 1 0 25424 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_279
timestamp 1663859327
transform 1 0 32592 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_283
timestamp 1663859327
transform 1 0 33040 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_286
timestamp 1663859327
transform 1 0 33376 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_350
timestamp 1663859327
transform 1 0 40544 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_354
timestamp 1663859327
transform 1 0 40992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_357
timestamp 1663859327
transform 1 0 41328 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_421
timestamp 1663859327
transform 1 0 48496 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_425
timestamp 1663859327
transform 1 0 48944 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_428
timestamp 1663859327
transform 1 0 49280 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_492
timestamp 1663859327
transform 1 0 56448 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_496
timestamp 1663859327
transform 1 0 56896 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_499
timestamp 1663859327
transform 1 0 57232 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_563
timestamp 1663859327
transform 1 0 64400 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_567
timestamp 1663859327
transform 1 0 64848 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_570
timestamp 1663859327
transform 1 0 65184 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_634
timestamp 1663859327
transform 1 0 72352 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_638
timestamp 1663859327
transform 1 0 72800 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_641
timestamp 1663859327
transform 1 0 73136 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_705
timestamp 1663859327
transform 1 0 80304 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_709
timestamp 1663859327
transform 1 0 80752 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_712
timestamp 1663859327
transform 1 0 81088 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_776
timestamp 1663859327
transform 1 0 88256 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_780
timestamp 1663859327
transform 1 0 88704 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_783
timestamp 1663859327
transform 1 0 89040 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_847
timestamp 1663859327
transform 1 0 96208 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_851
timestamp 1663859327
transform 1 0 96656 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_854
timestamp 1663859327
transform 1 0 96992 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_918
timestamp 1663859327
transform 1 0 104160 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_922
timestamp 1663859327
transform 1 0 104608 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_925
timestamp 1663859327
transform 1 0 104944 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_989
timestamp 1663859327
transform 1 0 112112 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_993
timestamp 1663859327
transform 1 0 112560 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_996
timestamp 1663859327
transform 1 0 112896 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_1028
timestamp 1663859327
transform 1 0 116480 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_1044
timestamp 1663859327
transform 1 0 118272 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_2
timestamp 1663859327
transform 1 0 1568 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_94_5
timestamp 1663859327
transform 1 0 1904 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_21
timestamp 1663859327
transform 1 0 3696 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_29
timestamp 1663859327
transform 1 0 4592 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_33
timestamp 1663859327
transform 1 0 5040 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_37
timestamp 1663859327
transform 1 0 5488 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_101
timestamp 1663859327
transform 1 0 12656 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_105
timestamp 1663859327
transform 1 0 13104 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_108
timestamp 1663859327
transform 1 0 13440 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_172
timestamp 1663859327
transform 1 0 20608 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_176
timestamp 1663859327
transform 1 0 21056 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_179
timestamp 1663859327
transform 1 0 21392 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_243
timestamp 1663859327
transform 1 0 28560 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_247
timestamp 1663859327
transform 1 0 29008 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_250
timestamp 1663859327
transform 1 0 29344 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_314
timestamp 1663859327
transform 1 0 36512 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_318
timestamp 1663859327
transform 1 0 36960 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_321
timestamp 1663859327
transform 1 0 37296 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_385
timestamp 1663859327
transform 1 0 44464 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_389
timestamp 1663859327
transform 1 0 44912 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_392
timestamp 1663859327
transform 1 0 45248 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_456
timestamp 1663859327
transform 1 0 52416 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_460
timestamp 1663859327
transform 1 0 52864 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_463
timestamp 1663859327
transform 1 0 53200 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_527
timestamp 1663859327
transform 1 0 60368 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_531
timestamp 1663859327
transform 1 0 60816 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_534
timestamp 1663859327
transform 1 0 61152 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_598
timestamp 1663859327
transform 1 0 68320 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_602
timestamp 1663859327
transform 1 0 68768 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_605
timestamp 1663859327
transform 1 0 69104 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_669
timestamp 1663859327
transform 1 0 76272 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_673
timestamp 1663859327
transform 1 0 76720 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_676
timestamp 1663859327
transform 1 0 77056 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_740
timestamp 1663859327
transform 1 0 84224 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_744
timestamp 1663859327
transform 1 0 84672 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_747
timestamp 1663859327
transform 1 0 85008 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_811
timestamp 1663859327
transform 1 0 92176 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_815
timestamp 1663859327
transform 1 0 92624 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_818
timestamp 1663859327
transform 1 0 92960 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_882
timestamp 1663859327
transform 1 0 100128 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_886
timestamp 1663859327
transform 1 0 100576 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_889
timestamp 1663859327
transform 1 0 100912 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_953
timestamp 1663859327
transform 1 0 108080 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_957
timestamp 1663859327
transform 1 0 108528 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_960
timestamp 1663859327
transform 1 0 108864 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_1024
timestamp 1663859327
transform 1 0 116032 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1028
timestamp 1663859327
transform 1 0 116480 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_1031
timestamp 1663859327
transform 1 0 116816 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1039
timestamp 1663859327
transform 1 0 117712 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_1044
timestamp 1663859327
transform 1 0 118272 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_2
timestamp 1663859327
transform 1 0 1568 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_95_9
timestamp 1663859327
transform 1 0 2352 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_95_41
timestamp 1663859327
transform 1 0 5936 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_57
timestamp 1663859327
transform 1 0 7728 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_65
timestamp 1663859327
transform 1 0 8624 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_69
timestamp 1663859327
transform 1 0 9072 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_73
timestamp 1663859327
transform 1 0 9520 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_137
timestamp 1663859327
transform 1 0 16688 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_141
timestamp 1663859327
transform 1 0 17136 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_144
timestamp 1663859327
transform 1 0 17472 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_208
timestamp 1663859327
transform 1 0 24640 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_212
timestamp 1663859327
transform 1 0 25088 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_215
timestamp 1663859327
transform 1 0 25424 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_279
timestamp 1663859327
transform 1 0 32592 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_283
timestamp 1663859327
transform 1 0 33040 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_286
timestamp 1663859327
transform 1 0 33376 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_350
timestamp 1663859327
transform 1 0 40544 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_354
timestamp 1663859327
transform 1 0 40992 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_357
timestamp 1663859327
transform 1 0 41328 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_421
timestamp 1663859327
transform 1 0 48496 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_425
timestamp 1663859327
transform 1 0 48944 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_428
timestamp 1663859327
transform 1 0 49280 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_492
timestamp 1663859327
transform 1 0 56448 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_496
timestamp 1663859327
transform 1 0 56896 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_499
timestamp 1663859327
transform 1 0 57232 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_563
timestamp 1663859327
transform 1 0 64400 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_567
timestamp 1663859327
transform 1 0 64848 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_570
timestamp 1663859327
transform 1 0 65184 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_634
timestamp 1663859327
transform 1 0 72352 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_638
timestamp 1663859327
transform 1 0 72800 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_641
timestamp 1663859327
transform 1 0 73136 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_705
timestamp 1663859327
transform 1 0 80304 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_709
timestamp 1663859327
transform 1 0 80752 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_712
timestamp 1663859327
transform 1 0 81088 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_776
timestamp 1663859327
transform 1 0 88256 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_780
timestamp 1663859327
transform 1 0 88704 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_783
timestamp 1663859327
transform 1 0 89040 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_847
timestamp 1663859327
transform 1 0 96208 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_851
timestamp 1663859327
transform 1 0 96656 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_854
timestamp 1663859327
transform 1 0 96992 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_918
timestamp 1663859327
transform 1 0 104160 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_922
timestamp 1663859327
transform 1 0 104608 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_925
timestamp 1663859327
transform 1 0 104944 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_989
timestamp 1663859327
transform 1 0 112112 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_993
timestamp 1663859327
transform 1 0 112560 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_95_996
timestamp 1663859327
transform 1 0 112896 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_95_1028
timestamp 1663859327
transform 1 0 116480 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_1044
timestamp 1663859327
transform 1 0 118272 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_96_2
timestamp 1663859327
transform 1 0 1568 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_34
timestamp 1663859327
transform 1 0 5152 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_37
timestamp 1663859327
transform 1 0 5488 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_101
timestamp 1663859327
transform 1 0 12656 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_105
timestamp 1663859327
transform 1 0 13104 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_108
timestamp 1663859327
transform 1 0 13440 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_172
timestamp 1663859327
transform 1 0 20608 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_176
timestamp 1663859327
transform 1 0 21056 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_179
timestamp 1663859327
transform 1 0 21392 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_243
timestamp 1663859327
transform 1 0 28560 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_247
timestamp 1663859327
transform 1 0 29008 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_250
timestamp 1663859327
transform 1 0 29344 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_314
timestamp 1663859327
transform 1 0 36512 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_318
timestamp 1663859327
transform 1 0 36960 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_321
timestamp 1663859327
transform 1 0 37296 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_385
timestamp 1663859327
transform 1 0 44464 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_389
timestamp 1663859327
transform 1 0 44912 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_392
timestamp 1663859327
transform 1 0 45248 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_456
timestamp 1663859327
transform 1 0 52416 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_460
timestamp 1663859327
transform 1 0 52864 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_463
timestamp 1663859327
transform 1 0 53200 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_527
timestamp 1663859327
transform 1 0 60368 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_531
timestamp 1663859327
transform 1 0 60816 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_534
timestamp 1663859327
transform 1 0 61152 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_598
timestamp 1663859327
transform 1 0 68320 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_602
timestamp 1663859327
transform 1 0 68768 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_605
timestamp 1663859327
transform 1 0 69104 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_669
timestamp 1663859327
transform 1 0 76272 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_673
timestamp 1663859327
transform 1 0 76720 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_676
timestamp 1663859327
transform 1 0 77056 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_740
timestamp 1663859327
transform 1 0 84224 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_744
timestamp 1663859327
transform 1 0 84672 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_747
timestamp 1663859327
transform 1 0 85008 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_811
timestamp 1663859327
transform 1 0 92176 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_815
timestamp 1663859327
transform 1 0 92624 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_818
timestamp 1663859327
transform 1 0 92960 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_882
timestamp 1663859327
transform 1 0 100128 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_886
timestamp 1663859327
transform 1 0 100576 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_889
timestamp 1663859327
transform 1 0 100912 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_953
timestamp 1663859327
transform 1 0 108080 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_957
timestamp 1663859327
transform 1 0 108528 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_960
timestamp 1663859327
transform 1 0 108864 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1024
timestamp 1663859327
transform 1 0 116032 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_1028
timestamp 1663859327
transform 1 0 116480 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_96_1031
timestamp 1663859327
transform 1 0 116816 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_1039
timestamp 1663859327
transform 1 0 117712 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_1043
timestamp 1663859327
transform 1 0 118160 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_2
timestamp 1663859327
transform 1 0 1568 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_66
timestamp 1663859327
transform 1 0 8736 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_70
timestamp 1663859327
transform 1 0 9184 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_73
timestamp 1663859327
transform 1 0 9520 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_137
timestamp 1663859327
transform 1 0 16688 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_141
timestamp 1663859327
transform 1 0 17136 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_144
timestamp 1663859327
transform 1 0 17472 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_208
timestamp 1663859327
transform 1 0 24640 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_212
timestamp 1663859327
transform 1 0 25088 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_215
timestamp 1663859327
transform 1 0 25424 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_279
timestamp 1663859327
transform 1 0 32592 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_283
timestamp 1663859327
transform 1 0 33040 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_286
timestamp 1663859327
transform 1 0 33376 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_350
timestamp 1663859327
transform 1 0 40544 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_354
timestamp 1663859327
transform 1 0 40992 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_357
timestamp 1663859327
transform 1 0 41328 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_421
timestamp 1663859327
transform 1 0 48496 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_425
timestamp 1663859327
transform 1 0 48944 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_428
timestamp 1663859327
transform 1 0 49280 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_492
timestamp 1663859327
transform 1 0 56448 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_496
timestamp 1663859327
transform 1 0 56896 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_499
timestamp 1663859327
transform 1 0 57232 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_563
timestamp 1663859327
transform 1 0 64400 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_567
timestamp 1663859327
transform 1 0 64848 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_570
timestamp 1663859327
transform 1 0 65184 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_634
timestamp 1663859327
transform 1 0 72352 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_638
timestamp 1663859327
transform 1 0 72800 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_641
timestamp 1663859327
transform 1 0 73136 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_705
timestamp 1663859327
transform 1 0 80304 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_709
timestamp 1663859327
transform 1 0 80752 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_712
timestamp 1663859327
transform 1 0 81088 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_776
timestamp 1663859327
transform 1 0 88256 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_780
timestamp 1663859327
transform 1 0 88704 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_783
timestamp 1663859327
transform 1 0 89040 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_847
timestamp 1663859327
transform 1 0 96208 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_851
timestamp 1663859327
transform 1 0 96656 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_854
timestamp 1663859327
transform 1 0 96992 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_918
timestamp 1663859327
transform 1 0 104160 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_922
timestamp 1663859327
transform 1 0 104608 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_925
timestamp 1663859327
transform 1 0 104944 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_989
timestamp 1663859327
transform 1 0 112112 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_993
timestamp 1663859327
transform 1 0 112560 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_97_996
timestamp 1663859327
transform 1 0 112896 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_97_1028
timestamp 1663859327
transform 1 0 116480 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_1036
timestamp 1663859327
transform 1 0 117376 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_1044
timestamp 1663859327
transform 1 0 118272 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_98_2
timestamp 1663859327
transform 1 0 1568 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_34
timestamp 1663859327
transform 1 0 5152 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_37
timestamp 1663859327
transform 1 0 5488 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_101
timestamp 1663859327
transform 1 0 12656 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_105
timestamp 1663859327
transform 1 0 13104 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_108
timestamp 1663859327
transform 1 0 13440 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_172
timestamp 1663859327
transform 1 0 20608 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_176
timestamp 1663859327
transform 1 0 21056 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_179
timestamp 1663859327
transform 1 0 21392 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_243
timestamp 1663859327
transform 1 0 28560 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_247
timestamp 1663859327
transform 1 0 29008 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_250
timestamp 1663859327
transform 1 0 29344 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_314
timestamp 1663859327
transform 1 0 36512 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_318
timestamp 1663859327
transform 1 0 36960 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_321
timestamp 1663859327
transform 1 0 37296 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_385
timestamp 1663859327
transform 1 0 44464 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_389
timestamp 1663859327
transform 1 0 44912 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_392
timestamp 1663859327
transform 1 0 45248 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_456
timestamp 1663859327
transform 1 0 52416 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_460
timestamp 1663859327
transform 1 0 52864 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_463
timestamp 1663859327
transform 1 0 53200 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_527
timestamp 1663859327
transform 1 0 60368 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_531
timestamp 1663859327
transform 1 0 60816 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_534
timestamp 1663859327
transform 1 0 61152 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_598
timestamp 1663859327
transform 1 0 68320 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_602
timestamp 1663859327
transform 1 0 68768 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_605
timestamp 1663859327
transform 1 0 69104 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_669
timestamp 1663859327
transform 1 0 76272 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_673
timestamp 1663859327
transform 1 0 76720 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_676
timestamp 1663859327
transform 1 0 77056 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_740
timestamp 1663859327
transform 1 0 84224 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_744
timestamp 1663859327
transform 1 0 84672 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_747
timestamp 1663859327
transform 1 0 85008 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_811
timestamp 1663859327
transform 1 0 92176 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_815
timestamp 1663859327
transform 1 0 92624 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_818
timestamp 1663859327
transform 1 0 92960 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_882
timestamp 1663859327
transform 1 0 100128 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_886
timestamp 1663859327
transform 1 0 100576 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_889
timestamp 1663859327
transform 1 0 100912 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_953
timestamp 1663859327
transform 1 0 108080 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_957
timestamp 1663859327
transform 1 0 108528 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_960
timestamp 1663859327
transform 1 0 108864 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1024
timestamp 1663859327
transform 1 0 116032 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_1028
timestamp 1663859327
transform 1 0 116480 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_98_1031
timestamp 1663859327
transform 1 0 116816 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_1039
timestamp 1663859327
transform 1 0 117712 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_1043
timestamp 1663859327
transform 1 0 118160 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_2
timestamp 1663859327
transform 1 0 1568 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_66
timestamp 1663859327
transform 1 0 8736 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_70
timestamp 1663859327
transform 1 0 9184 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_73
timestamp 1663859327
transform 1 0 9520 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_137
timestamp 1663859327
transform 1 0 16688 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_141
timestamp 1663859327
transform 1 0 17136 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_144
timestamp 1663859327
transform 1 0 17472 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_208
timestamp 1663859327
transform 1 0 24640 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_212
timestamp 1663859327
transform 1 0 25088 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_215
timestamp 1663859327
transform 1 0 25424 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_279
timestamp 1663859327
transform 1 0 32592 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_283
timestamp 1663859327
transform 1 0 33040 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_286
timestamp 1663859327
transform 1 0 33376 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_350
timestamp 1663859327
transform 1 0 40544 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_354
timestamp 1663859327
transform 1 0 40992 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_357
timestamp 1663859327
transform 1 0 41328 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_421
timestamp 1663859327
transform 1 0 48496 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_425
timestamp 1663859327
transform 1 0 48944 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_428
timestamp 1663859327
transform 1 0 49280 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_492
timestamp 1663859327
transform 1 0 56448 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_496
timestamp 1663859327
transform 1 0 56896 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_499
timestamp 1663859327
transform 1 0 57232 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_563
timestamp 1663859327
transform 1 0 64400 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_567
timestamp 1663859327
transform 1 0 64848 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_570
timestamp 1663859327
transform 1 0 65184 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_634
timestamp 1663859327
transform 1 0 72352 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_638
timestamp 1663859327
transform 1 0 72800 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_641
timestamp 1663859327
transform 1 0 73136 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_705
timestamp 1663859327
transform 1 0 80304 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_709
timestamp 1663859327
transform 1 0 80752 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_712
timestamp 1663859327
transform 1 0 81088 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_776
timestamp 1663859327
transform 1 0 88256 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_780
timestamp 1663859327
transform 1 0 88704 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_783
timestamp 1663859327
transform 1 0 89040 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_847
timestamp 1663859327
transform 1 0 96208 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_851
timestamp 1663859327
transform 1 0 96656 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_854
timestamp 1663859327
transform 1 0 96992 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_918
timestamp 1663859327
transform 1 0 104160 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_922
timestamp 1663859327
transform 1 0 104608 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_925
timestamp 1663859327
transform 1 0 104944 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_989
timestamp 1663859327
transform 1 0 112112 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_993
timestamp 1663859327
transform 1 0 112560 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_99_996
timestamp 1663859327
transform 1 0 112896 0 -1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_99_1028
timestamp 1663859327
transform 1 0 116480 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_1044
timestamp 1663859327
transform 1 0 118272 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_100_2
timestamp 1663859327
transform 1 0 1568 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_34
timestamp 1663859327
transform 1 0 5152 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_37
timestamp 1663859327
transform 1 0 5488 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_101
timestamp 1663859327
transform 1 0 12656 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_105
timestamp 1663859327
transform 1 0 13104 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_108
timestamp 1663859327
transform 1 0 13440 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_172
timestamp 1663859327
transform 1 0 20608 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_176
timestamp 1663859327
transform 1 0 21056 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_179
timestamp 1663859327
transform 1 0 21392 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_243
timestamp 1663859327
transform 1 0 28560 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_247
timestamp 1663859327
transform 1 0 29008 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_250
timestamp 1663859327
transform 1 0 29344 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_314
timestamp 1663859327
transform 1 0 36512 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_318
timestamp 1663859327
transform 1 0 36960 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_321
timestamp 1663859327
transform 1 0 37296 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_385
timestamp 1663859327
transform 1 0 44464 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_389
timestamp 1663859327
transform 1 0 44912 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_392
timestamp 1663859327
transform 1 0 45248 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_456
timestamp 1663859327
transform 1 0 52416 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_460
timestamp 1663859327
transform 1 0 52864 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_463
timestamp 1663859327
transform 1 0 53200 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_527
timestamp 1663859327
transform 1 0 60368 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_531
timestamp 1663859327
transform 1 0 60816 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_534
timestamp 1663859327
transform 1 0 61152 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_598
timestamp 1663859327
transform 1 0 68320 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_602
timestamp 1663859327
transform 1 0 68768 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_605
timestamp 1663859327
transform 1 0 69104 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_669
timestamp 1663859327
transform 1 0 76272 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_673
timestamp 1663859327
transform 1 0 76720 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_676
timestamp 1663859327
transform 1 0 77056 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_740
timestamp 1663859327
transform 1 0 84224 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_744
timestamp 1663859327
transform 1 0 84672 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_747
timestamp 1663859327
transform 1 0 85008 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_811
timestamp 1663859327
transform 1 0 92176 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_815
timestamp 1663859327
transform 1 0 92624 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_818
timestamp 1663859327
transform 1 0 92960 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_882
timestamp 1663859327
transform 1 0 100128 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_886
timestamp 1663859327
transform 1 0 100576 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_889
timestamp 1663859327
transform 1 0 100912 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_953
timestamp 1663859327
transform 1 0 108080 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_957
timestamp 1663859327
transform 1 0 108528 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_960
timestamp 1663859327
transform 1 0 108864 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1024
timestamp 1663859327
transform 1 0 116032 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_1028
timestamp 1663859327
transform 1 0 116480 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_1031
timestamp 1663859327
transform 1 0 116816 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_1039
timestamp 1663859327
transform 1 0 117712 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_1043
timestamp 1663859327
transform 1 0 118160 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_2
timestamp 1663859327
transform 1 0 1568 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_66
timestamp 1663859327
transform 1 0 8736 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_70
timestamp 1663859327
transform 1 0 9184 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_73
timestamp 1663859327
transform 1 0 9520 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_137
timestamp 1663859327
transform 1 0 16688 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_141
timestamp 1663859327
transform 1 0 17136 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_144
timestamp 1663859327
transform 1 0 17472 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_208
timestamp 1663859327
transform 1 0 24640 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_212
timestamp 1663859327
transform 1 0 25088 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_215
timestamp 1663859327
transform 1 0 25424 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_279
timestamp 1663859327
transform 1 0 32592 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_283
timestamp 1663859327
transform 1 0 33040 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_286
timestamp 1663859327
transform 1 0 33376 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_350
timestamp 1663859327
transform 1 0 40544 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_354
timestamp 1663859327
transform 1 0 40992 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_357
timestamp 1663859327
transform 1 0 41328 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_421
timestamp 1663859327
transform 1 0 48496 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_425
timestamp 1663859327
transform 1 0 48944 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_428
timestamp 1663859327
transform 1 0 49280 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_492
timestamp 1663859327
transform 1 0 56448 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_496
timestamp 1663859327
transform 1 0 56896 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_499
timestamp 1663859327
transform 1 0 57232 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_563
timestamp 1663859327
transform 1 0 64400 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_567
timestamp 1663859327
transform 1 0 64848 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_570
timestamp 1663859327
transform 1 0 65184 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_634
timestamp 1663859327
transform 1 0 72352 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_638
timestamp 1663859327
transform 1 0 72800 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_641
timestamp 1663859327
transform 1 0 73136 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_705
timestamp 1663859327
transform 1 0 80304 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_709
timestamp 1663859327
transform 1 0 80752 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_712
timestamp 1663859327
transform 1 0 81088 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_776
timestamp 1663859327
transform 1 0 88256 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_780
timestamp 1663859327
transform 1 0 88704 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_783
timestamp 1663859327
transform 1 0 89040 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_847
timestamp 1663859327
transform 1 0 96208 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_851
timestamp 1663859327
transform 1 0 96656 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_854
timestamp 1663859327
transform 1 0 96992 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_918
timestamp 1663859327
transform 1 0 104160 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_922
timestamp 1663859327
transform 1 0 104608 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_925
timestamp 1663859327
transform 1 0 104944 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_989
timestamp 1663859327
transform 1 0 112112 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_993
timestamp 1663859327
transform 1 0 112560 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_101_996
timestamp 1663859327
transform 1 0 112896 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_1028
timestamp 1663859327
transform 1 0 116480 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_1036
timestamp 1663859327
transform 1 0 117376 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_1044
timestamp 1663859327
transform 1 0 118272 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_2
timestamp 1663859327
transform 1 0 1568 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_7
timestamp 1663859327
transform 1 0 2128 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_13
timestamp 1663859327
transform 1 0 2800 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_29
timestamp 1663859327
transform 1 0 4592 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_33
timestamp 1663859327
transform 1 0 5040 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_37
timestamp 1663859327
transform 1 0 5488 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_101
timestamp 1663859327
transform 1 0 12656 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_105
timestamp 1663859327
transform 1 0 13104 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_108
timestamp 1663859327
transform 1 0 13440 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_172
timestamp 1663859327
transform 1 0 20608 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_176
timestamp 1663859327
transform 1 0 21056 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_179
timestamp 1663859327
transform 1 0 21392 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_243
timestamp 1663859327
transform 1 0 28560 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_247
timestamp 1663859327
transform 1 0 29008 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_250
timestamp 1663859327
transform 1 0 29344 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_314
timestamp 1663859327
transform 1 0 36512 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_318
timestamp 1663859327
transform 1 0 36960 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_321
timestamp 1663859327
transform 1 0 37296 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_385
timestamp 1663859327
transform 1 0 44464 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_389
timestamp 1663859327
transform 1 0 44912 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_392
timestamp 1663859327
transform 1 0 45248 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_456
timestamp 1663859327
transform 1 0 52416 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_460
timestamp 1663859327
transform 1 0 52864 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_463
timestamp 1663859327
transform 1 0 53200 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_527
timestamp 1663859327
transform 1 0 60368 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_531
timestamp 1663859327
transform 1 0 60816 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_534
timestamp 1663859327
transform 1 0 61152 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_598
timestamp 1663859327
transform 1 0 68320 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_602
timestamp 1663859327
transform 1 0 68768 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_605
timestamp 1663859327
transform 1 0 69104 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_669
timestamp 1663859327
transform 1 0 76272 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_673
timestamp 1663859327
transform 1 0 76720 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_676
timestamp 1663859327
transform 1 0 77056 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_740
timestamp 1663859327
transform 1 0 84224 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_744
timestamp 1663859327
transform 1 0 84672 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_747
timestamp 1663859327
transform 1 0 85008 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_811
timestamp 1663859327
transform 1 0 92176 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_815
timestamp 1663859327
transform 1 0 92624 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_818
timestamp 1663859327
transform 1 0 92960 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_882
timestamp 1663859327
transform 1 0 100128 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_886
timestamp 1663859327
transform 1 0 100576 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_889
timestamp 1663859327
transform 1 0 100912 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_953
timestamp 1663859327
transform 1 0 108080 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_957
timestamp 1663859327
transform 1 0 108528 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_960
timestamp 1663859327
transform 1 0 108864 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1024
timestamp 1663859327
transform 1 0 116032 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_1028
timestamp 1663859327
transform 1 0 116480 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_102_1031
timestamp 1663859327
transform 1 0 116816 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_1039
timestamp 1663859327
transform 1 0 117712 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_1043
timestamp 1663859327
transform 1 0 118160 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_2
timestamp 1663859327
transform 1 0 1568 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_66
timestamp 1663859327
transform 1 0 8736 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_70
timestamp 1663859327
transform 1 0 9184 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_73
timestamp 1663859327
transform 1 0 9520 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_137
timestamp 1663859327
transform 1 0 16688 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_141
timestamp 1663859327
transform 1 0 17136 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_144
timestamp 1663859327
transform 1 0 17472 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_208
timestamp 1663859327
transform 1 0 24640 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_212
timestamp 1663859327
transform 1 0 25088 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_215
timestamp 1663859327
transform 1 0 25424 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_279
timestamp 1663859327
transform 1 0 32592 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_283
timestamp 1663859327
transform 1 0 33040 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_286
timestamp 1663859327
transform 1 0 33376 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_350
timestamp 1663859327
transform 1 0 40544 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_354
timestamp 1663859327
transform 1 0 40992 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_357
timestamp 1663859327
transform 1 0 41328 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_421
timestamp 1663859327
transform 1 0 48496 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_425
timestamp 1663859327
transform 1 0 48944 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_428
timestamp 1663859327
transform 1 0 49280 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_492
timestamp 1663859327
transform 1 0 56448 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_496
timestamp 1663859327
transform 1 0 56896 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_499
timestamp 1663859327
transform 1 0 57232 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_563
timestamp 1663859327
transform 1 0 64400 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_567
timestamp 1663859327
transform 1 0 64848 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_570
timestamp 1663859327
transform 1 0 65184 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_634
timestamp 1663859327
transform 1 0 72352 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_638
timestamp 1663859327
transform 1 0 72800 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_641
timestamp 1663859327
transform 1 0 73136 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_705
timestamp 1663859327
transform 1 0 80304 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_709
timestamp 1663859327
transform 1 0 80752 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_712
timestamp 1663859327
transform 1 0 81088 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_776
timestamp 1663859327
transform 1 0 88256 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_780
timestamp 1663859327
transform 1 0 88704 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_783
timestamp 1663859327
transform 1 0 89040 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_847
timestamp 1663859327
transform 1 0 96208 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_851
timestamp 1663859327
transform 1 0 96656 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_854
timestamp 1663859327
transform 1 0 96992 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_918
timestamp 1663859327
transform 1 0 104160 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_922
timestamp 1663859327
transform 1 0 104608 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_925
timestamp 1663859327
transform 1 0 104944 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_989
timestamp 1663859327
transform 1 0 112112 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_993
timestamp 1663859327
transform 1 0 112560 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_103_996
timestamp 1663859327
transform 1 0 112896 0 -1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_103_1028
timestamp 1663859327
transform 1 0 116480 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_1036
timestamp 1663859327
transform 1 0 117376 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_1044
timestamp 1663859327
transform 1 0 118272 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_2
timestamp 1663859327
transform 1 0 1568 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_17
timestamp 1663859327
transform 1 0 3248 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_21
timestamp 1663859327
transform 1 0 3696 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_29
timestamp 1663859327
transform 1 0 4592 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_33
timestamp 1663859327
transform 1 0 5040 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_37
timestamp 1663859327
transform 1 0 5488 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_101
timestamp 1663859327
transform 1 0 12656 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_105
timestamp 1663859327
transform 1 0 13104 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_108
timestamp 1663859327
transform 1 0 13440 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_172
timestamp 1663859327
transform 1 0 20608 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_176
timestamp 1663859327
transform 1 0 21056 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_179
timestamp 1663859327
transform 1 0 21392 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_243
timestamp 1663859327
transform 1 0 28560 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_247
timestamp 1663859327
transform 1 0 29008 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_250
timestamp 1663859327
transform 1 0 29344 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_314
timestamp 1663859327
transform 1 0 36512 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_318
timestamp 1663859327
transform 1 0 36960 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_321
timestamp 1663859327
transform 1 0 37296 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_385
timestamp 1663859327
transform 1 0 44464 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_389
timestamp 1663859327
transform 1 0 44912 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_392
timestamp 1663859327
transform 1 0 45248 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_456
timestamp 1663859327
transform 1 0 52416 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_460
timestamp 1663859327
transform 1 0 52864 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_463
timestamp 1663859327
transform 1 0 53200 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_527
timestamp 1663859327
transform 1 0 60368 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_531
timestamp 1663859327
transform 1 0 60816 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_534
timestamp 1663859327
transform 1 0 61152 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_598
timestamp 1663859327
transform 1 0 68320 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_602
timestamp 1663859327
transform 1 0 68768 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_605
timestamp 1663859327
transform 1 0 69104 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_669
timestamp 1663859327
transform 1 0 76272 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_673
timestamp 1663859327
transform 1 0 76720 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_676
timestamp 1663859327
transform 1 0 77056 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_740
timestamp 1663859327
transform 1 0 84224 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_744
timestamp 1663859327
transform 1 0 84672 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_747
timestamp 1663859327
transform 1 0 85008 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_811
timestamp 1663859327
transform 1 0 92176 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_815
timestamp 1663859327
transform 1 0 92624 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_818
timestamp 1663859327
transform 1 0 92960 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_882
timestamp 1663859327
transform 1 0 100128 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_886
timestamp 1663859327
transform 1 0 100576 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_889
timestamp 1663859327
transform 1 0 100912 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_953
timestamp 1663859327
transform 1 0 108080 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_957
timestamp 1663859327
transform 1 0 108528 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_960
timestamp 1663859327
transform 1 0 108864 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1024
timestamp 1663859327
transform 1 0 116032 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_1028
timestamp 1663859327
transform 1 0 116480 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_1031
timestamp 1663859327
transform 1 0 116816 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_1039
timestamp 1663859327
transform 1 0 117712 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_1043
timestamp 1663859327
transform 1 0 118160 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_2
timestamp 1663859327
transform 1 0 1568 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_66
timestamp 1663859327
transform 1 0 8736 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_70
timestamp 1663859327
transform 1 0 9184 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_73
timestamp 1663859327
transform 1 0 9520 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_137
timestamp 1663859327
transform 1 0 16688 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_141
timestamp 1663859327
transform 1 0 17136 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_144
timestamp 1663859327
transform 1 0 17472 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_208
timestamp 1663859327
transform 1 0 24640 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_212
timestamp 1663859327
transform 1 0 25088 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_215
timestamp 1663859327
transform 1 0 25424 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_279
timestamp 1663859327
transform 1 0 32592 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_283
timestamp 1663859327
transform 1 0 33040 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_286
timestamp 1663859327
transform 1 0 33376 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_350
timestamp 1663859327
transform 1 0 40544 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_354
timestamp 1663859327
transform 1 0 40992 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_357
timestamp 1663859327
transform 1 0 41328 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_421
timestamp 1663859327
transform 1 0 48496 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_425
timestamp 1663859327
transform 1 0 48944 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_428
timestamp 1663859327
transform 1 0 49280 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_492
timestamp 1663859327
transform 1 0 56448 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_496
timestamp 1663859327
transform 1 0 56896 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_499
timestamp 1663859327
transform 1 0 57232 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_563
timestamp 1663859327
transform 1 0 64400 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_567
timestamp 1663859327
transform 1 0 64848 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_570
timestamp 1663859327
transform 1 0 65184 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_634
timestamp 1663859327
transform 1 0 72352 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_638
timestamp 1663859327
transform 1 0 72800 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_641
timestamp 1663859327
transform 1 0 73136 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_705
timestamp 1663859327
transform 1 0 80304 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_709
timestamp 1663859327
transform 1 0 80752 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_712
timestamp 1663859327
transform 1 0 81088 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_776
timestamp 1663859327
transform 1 0 88256 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_780
timestamp 1663859327
transform 1 0 88704 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_783
timestamp 1663859327
transform 1 0 89040 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_847
timestamp 1663859327
transform 1 0 96208 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_851
timestamp 1663859327
transform 1 0 96656 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_854
timestamp 1663859327
transform 1 0 96992 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_918
timestamp 1663859327
transform 1 0 104160 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_922
timestamp 1663859327
transform 1 0 104608 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_925
timestamp 1663859327
transform 1 0 104944 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_989
timestamp 1663859327
transform 1 0 112112 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_993
timestamp 1663859327
transform 1 0 112560 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_105_996
timestamp 1663859327
transform 1 0 112896 0 -1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_105_1028
timestamp 1663859327
transform 1 0 116480 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_1044
timestamp 1663859327
transform 1 0 118272 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_106_2
timestamp 1663859327
transform 1 0 1568 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_34
timestamp 1663859327
transform 1 0 5152 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_37
timestamp 1663859327
transform 1 0 5488 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_101
timestamp 1663859327
transform 1 0 12656 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_105
timestamp 1663859327
transform 1 0 13104 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_108
timestamp 1663859327
transform 1 0 13440 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_172
timestamp 1663859327
transform 1 0 20608 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_176
timestamp 1663859327
transform 1 0 21056 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_179
timestamp 1663859327
transform 1 0 21392 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_243
timestamp 1663859327
transform 1 0 28560 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_247
timestamp 1663859327
transform 1 0 29008 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_250
timestamp 1663859327
transform 1 0 29344 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_314
timestamp 1663859327
transform 1 0 36512 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_318
timestamp 1663859327
transform 1 0 36960 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_321
timestamp 1663859327
transform 1 0 37296 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_385
timestamp 1663859327
transform 1 0 44464 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_389
timestamp 1663859327
transform 1 0 44912 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_392
timestamp 1663859327
transform 1 0 45248 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_456
timestamp 1663859327
transform 1 0 52416 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_460
timestamp 1663859327
transform 1 0 52864 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_463
timestamp 1663859327
transform 1 0 53200 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_527
timestamp 1663859327
transform 1 0 60368 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_531
timestamp 1663859327
transform 1 0 60816 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_534
timestamp 1663859327
transform 1 0 61152 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_598
timestamp 1663859327
transform 1 0 68320 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_602
timestamp 1663859327
transform 1 0 68768 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_605
timestamp 1663859327
transform 1 0 69104 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_669
timestamp 1663859327
transform 1 0 76272 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_673
timestamp 1663859327
transform 1 0 76720 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_676
timestamp 1663859327
transform 1 0 77056 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_740
timestamp 1663859327
transform 1 0 84224 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_744
timestamp 1663859327
transform 1 0 84672 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_747
timestamp 1663859327
transform 1 0 85008 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_811
timestamp 1663859327
transform 1 0 92176 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_815
timestamp 1663859327
transform 1 0 92624 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_818
timestamp 1663859327
transform 1 0 92960 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_882
timestamp 1663859327
transform 1 0 100128 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_886
timestamp 1663859327
transform 1 0 100576 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_889
timestamp 1663859327
transform 1 0 100912 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_953
timestamp 1663859327
transform 1 0 108080 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_957
timestamp 1663859327
transform 1 0 108528 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_960
timestamp 1663859327
transform 1 0 108864 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1024
timestamp 1663859327
transform 1 0 116032 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_1028
timestamp 1663859327
transform 1 0 116480 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_1031
timestamp 1663859327
transform 1 0 116816 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_1039
timestamp 1663859327
transform 1 0 117712 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_1043
timestamp 1663859327
transform 1 0 118160 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_2
timestamp 1663859327
transform 1 0 1568 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_66
timestamp 1663859327
transform 1 0 8736 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_70
timestamp 1663859327
transform 1 0 9184 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_73
timestamp 1663859327
transform 1 0 9520 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_137
timestamp 1663859327
transform 1 0 16688 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_141
timestamp 1663859327
transform 1 0 17136 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_144
timestamp 1663859327
transform 1 0 17472 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_208
timestamp 1663859327
transform 1 0 24640 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_212
timestamp 1663859327
transform 1 0 25088 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_215
timestamp 1663859327
transform 1 0 25424 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_279
timestamp 1663859327
transform 1 0 32592 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_283
timestamp 1663859327
transform 1 0 33040 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_286
timestamp 1663859327
transform 1 0 33376 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_350
timestamp 1663859327
transform 1 0 40544 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_354
timestamp 1663859327
transform 1 0 40992 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_357
timestamp 1663859327
transform 1 0 41328 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_421
timestamp 1663859327
transform 1 0 48496 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_425
timestamp 1663859327
transform 1 0 48944 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_428
timestamp 1663859327
transform 1 0 49280 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_492
timestamp 1663859327
transform 1 0 56448 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_496
timestamp 1663859327
transform 1 0 56896 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_499
timestamp 1663859327
transform 1 0 57232 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_563
timestamp 1663859327
transform 1 0 64400 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_567
timestamp 1663859327
transform 1 0 64848 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_570
timestamp 1663859327
transform 1 0 65184 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_634
timestamp 1663859327
transform 1 0 72352 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_638
timestamp 1663859327
transform 1 0 72800 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_641
timestamp 1663859327
transform 1 0 73136 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_705
timestamp 1663859327
transform 1 0 80304 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_709
timestamp 1663859327
transform 1 0 80752 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_712
timestamp 1663859327
transform 1 0 81088 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_776
timestamp 1663859327
transform 1 0 88256 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_780
timestamp 1663859327
transform 1 0 88704 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_783
timestamp 1663859327
transform 1 0 89040 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_847
timestamp 1663859327
transform 1 0 96208 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_851
timestamp 1663859327
transform 1 0 96656 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_854
timestamp 1663859327
transform 1 0 96992 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_918
timestamp 1663859327
transform 1 0 104160 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_922
timestamp 1663859327
transform 1 0 104608 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_925
timestamp 1663859327
transform 1 0 104944 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_989
timestamp 1663859327
transform 1 0 112112 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_993
timestamp 1663859327
transform 1 0 112560 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_107_996
timestamp 1663859327
transform 1 0 112896 0 -1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_107_1028
timestamp 1663859327
transform 1 0 116480 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_1044
timestamp 1663859327
transform 1 0 118272 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_108_2
timestamp 1663859327
transform 1 0 1568 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_34
timestamp 1663859327
transform 1 0 5152 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_37
timestamp 1663859327
transform 1 0 5488 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_101
timestamp 1663859327
transform 1 0 12656 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_105
timestamp 1663859327
transform 1 0 13104 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_108
timestamp 1663859327
transform 1 0 13440 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_172
timestamp 1663859327
transform 1 0 20608 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_176
timestamp 1663859327
transform 1 0 21056 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_179
timestamp 1663859327
transform 1 0 21392 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_243
timestamp 1663859327
transform 1 0 28560 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_247
timestamp 1663859327
transform 1 0 29008 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_250
timestamp 1663859327
transform 1 0 29344 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_314
timestamp 1663859327
transform 1 0 36512 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_318
timestamp 1663859327
transform 1 0 36960 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_321
timestamp 1663859327
transform 1 0 37296 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_385
timestamp 1663859327
transform 1 0 44464 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_389
timestamp 1663859327
transform 1 0 44912 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_392
timestamp 1663859327
transform 1 0 45248 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_456
timestamp 1663859327
transform 1 0 52416 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_460
timestamp 1663859327
transform 1 0 52864 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_463
timestamp 1663859327
transform 1 0 53200 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_527
timestamp 1663859327
transform 1 0 60368 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_531
timestamp 1663859327
transform 1 0 60816 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_534
timestamp 1663859327
transform 1 0 61152 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_598
timestamp 1663859327
transform 1 0 68320 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_602
timestamp 1663859327
transform 1 0 68768 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_605
timestamp 1663859327
transform 1 0 69104 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_669
timestamp 1663859327
transform 1 0 76272 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_673
timestamp 1663859327
transform 1 0 76720 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_676
timestamp 1663859327
transform 1 0 77056 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_740
timestamp 1663859327
transform 1 0 84224 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_744
timestamp 1663859327
transform 1 0 84672 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_747
timestamp 1663859327
transform 1 0 85008 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_811
timestamp 1663859327
transform 1 0 92176 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_815
timestamp 1663859327
transform 1 0 92624 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_818
timestamp 1663859327
transform 1 0 92960 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_882
timestamp 1663859327
transform 1 0 100128 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_886
timestamp 1663859327
transform 1 0 100576 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_889
timestamp 1663859327
transform 1 0 100912 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_953
timestamp 1663859327
transform 1 0 108080 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_957
timestamp 1663859327
transform 1 0 108528 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_960
timestamp 1663859327
transform 1 0 108864 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_1024
timestamp 1663859327
transform 1 0 116032 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1028
timestamp 1663859327
transform 1 0 116480 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_108_1031
timestamp 1663859327
transform 1 0 116816 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1039
timestamp 1663859327
transform 1 0 117712 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_1044
timestamp 1663859327
transform 1 0 118272 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_2
timestamp 1663859327
transform 1 0 1568 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_66
timestamp 1663859327
transform 1 0 8736 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_70
timestamp 1663859327
transform 1 0 9184 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_73
timestamp 1663859327
transform 1 0 9520 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_137
timestamp 1663859327
transform 1 0 16688 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_141
timestamp 1663859327
transform 1 0 17136 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_144
timestamp 1663859327
transform 1 0 17472 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_208
timestamp 1663859327
transform 1 0 24640 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_212
timestamp 1663859327
transform 1 0 25088 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_215
timestamp 1663859327
transform 1 0 25424 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_279
timestamp 1663859327
transform 1 0 32592 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_283
timestamp 1663859327
transform 1 0 33040 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_286
timestamp 1663859327
transform 1 0 33376 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_350
timestamp 1663859327
transform 1 0 40544 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_354
timestamp 1663859327
transform 1 0 40992 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_357
timestamp 1663859327
transform 1 0 41328 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_421
timestamp 1663859327
transform 1 0 48496 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_425
timestamp 1663859327
transform 1 0 48944 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_428
timestamp 1663859327
transform 1 0 49280 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_492
timestamp 1663859327
transform 1 0 56448 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_496
timestamp 1663859327
transform 1 0 56896 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_499
timestamp 1663859327
transform 1 0 57232 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_563
timestamp 1663859327
transform 1 0 64400 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_567
timestamp 1663859327
transform 1 0 64848 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_570
timestamp 1663859327
transform 1 0 65184 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_634
timestamp 1663859327
transform 1 0 72352 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_638
timestamp 1663859327
transform 1 0 72800 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_641
timestamp 1663859327
transform 1 0 73136 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_705
timestamp 1663859327
transform 1 0 80304 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_709
timestamp 1663859327
transform 1 0 80752 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_712
timestamp 1663859327
transform 1 0 81088 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_776
timestamp 1663859327
transform 1 0 88256 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_780
timestamp 1663859327
transform 1 0 88704 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_783
timestamp 1663859327
transform 1 0 89040 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_847
timestamp 1663859327
transform 1 0 96208 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_851
timestamp 1663859327
transform 1 0 96656 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_854
timestamp 1663859327
transform 1 0 96992 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_918
timestamp 1663859327
transform 1 0 104160 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_922
timestamp 1663859327
transform 1 0 104608 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_925
timestamp 1663859327
transform 1 0 104944 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_989
timestamp 1663859327
transform 1 0 112112 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_993
timestamp 1663859327
transform 1 0 112560 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_109_996
timestamp 1663859327
transform 1 0 112896 0 -1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_1028
timestamp 1663859327
transform 1 0 116480 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_1044
timestamp 1663859327
transform 1 0 118272 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_2
timestamp 1663859327
transform 1 0 1568 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_110_5
timestamp 1663859327
transform 1 0 1904 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_110_21
timestamp 1663859327
transform 1 0 3696 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_29
timestamp 1663859327
transform 1 0 4592 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_33
timestamp 1663859327
transform 1 0 5040 0 1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_37
timestamp 1663859327
transform 1 0 5488 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_101
timestamp 1663859327
transform 1 0 12656 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_105
timestamp 1663859327
transform 1 0 13104 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_108
timestamp 1663859327
transform 1 0 13440 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_172
timestamp 1663859327
transform 1 0 20608 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_176
timestamp 1663859327
transform 1 0 21056 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_179
timestamp 1663859327
transform 1 0 21392 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_243
timestamp 1663859327
transform 1 0 28560 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_247
timestamp 1663859327
transform 1 0 29008 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_250
timestamp 1663859327
transform 1 0 29344 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_314
timestamp 1663859327
transform 1 0 36512 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_318
timestamp 1663859327
transform 1 0 36960 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_321
timestamp 1663859327
transform 1 0 37296 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_385
timestamp 1663859327
transform 1 0 44464 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_389
timestamp 1663859327
transform 1 0 44912 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_392
timestamp 1663859327
transform 1 0 45248 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_456
timestamp 1663859327
transform 1 0 52416 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_460
timestamp 1663859327
transform 1 0 52864 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_463
timestamp 1663859327
transform 1 0 53200 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_527
timestamp 1663859327
transform 1 0 60368 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_531
timestamp 1663859327
transform 1 0 60816 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_534
timestamp 1663859327
transform 1 0 61152 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_598
timestamp 1663859327
transform 1 0 68320 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_602
timestamp 1663859327
transform 1 0 68768 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_605
timestamp 1663859327
transform 1 0 69104 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_669
timestamp 1663859327
transform 1 0 76272 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_673
timestamp 1663859327
transform 1 0 76720 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_676
timestamp 1663859327
transform 1 0 77056 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_740
timestamp 1663859327
transform 1 0 84224 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_744
timestamp 1663859327
transform 1 0 84672 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_747
timestamp 1663859327
transform 1 0 85008 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_811
timestamp 1663859327
transform 1 0 92176 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_815
timestamp 1663859327
transform 1 0 92624 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_818
timestamp 1663859327
transform 1 0 92960 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_882
timestamp 1663859327
transform 1 0 100128 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_886
timestamp 1663859327
transform 1 0 100576 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_889
timestamp 1663859327
transform 1 0 100912 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_953
timestamp 1663859327
transform 1 0 108080 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_957
timestamp 1663859327
transform 1 0 108528 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_960
timestamp 1663859327
transform 1 0 108864 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1024
timestamp 1663859327
transform 1 0 116032 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_1028
timestamp 1663859327
transform 1 0 116480 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_110_1031
timestamp 1663859327
transform 1 0 116816 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_1039
timestamp 1663859327
transform 1 0 117712 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_1043
timestamp 1663859327
transform 1 0 118160 0 1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_2
timestamp 1663859327
transform 1 0 1568 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_111_9
timestamp 1663859327
transform 1 0 2352 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_111_41
timestamp 1663859327
transform 1 0 5936 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_111_57
timestamp 1663859327
transform 1 0 7728 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_65
timestamp 1663859327
transform 1 0 8624 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_111_69
timestamp 1663859327
transform 1 0 9072 0 -1 90944
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_73
timestamp 1663859327
transform 1 0 9520 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_137
timestamp 1663859327
transform 1 0 16688 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_141
timestamp 1663859327
transform 1 0 17136 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_144
timestamp 1663859327
transform 1 0 17472 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_208
timestamp 1663859327
transform 1 0 24640 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_212
timestamp 1663859327
transform 1 0 25088 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_215
timestamp 1663859327
transform 1 0 25424 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_279
timestamp 1663859327
transform 1 0 32592 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_283
timestamp 1663859327
transform 1 0 33040 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_286
timestamp 1663859327
transform 1 0 33376 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_350
timestamp 1663859327
transform 1 0 40544 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_354
timestamp 1663859327
transform 1 0 40992 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_357
timestamp 1663859327
transform 1 0 41328 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_421
timestamp 1663859327
transform 1 0 48496 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_425
timestamp 1663859327
transform 1 0 48944 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_428
timestamp 1663859327
transform 1 0 49280 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_492
timestamp 1663859327
transform 1 0 56448 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_496
timestamp 1663859327
transform 1 0 56896 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_499
timestamp 1663859327
transform 1 0 57232 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_563
timestamp 1663859327
transform 1 0 64400 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_567
timestamp 1663859327
transform 1 0 64848 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_570
timestamp 1663859327
transform 1 0 65184 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_634
timestamp 1663859327
transform 1 0 72352 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_638
timestamp 1663859327
transform 1 0 72800 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_641
timestamp 1663859327
transform 1 0 73136 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_705
timestamp 1663859327
transform 1 0 80304 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_709
timestamp 1663859327
transform 1 0 80752 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_712
timestamp 1663859327
transform 1 0 81088 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_776
timestamp 1663859327
transform 1 0 88256 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_780
timestamp 1663859327
transform 1 0 88704 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_783
timestamp 1663859327
transform 1 0 89040 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_847
timestamp 1663859327
transform 1 0 96208 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_851
timestamp 1663859327
transform 1 0 96656 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_854
timestamp 1663859327
transform 1 0 96992 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_918
timestamp 1663859327
transform 1 0 104160 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_922
timestamp 1663859327
transform 1 0 104608 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_925
timestamp 1663859327
transform 1 0 104944 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_989
timestamp 1663859327
transform 1 0 112112 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_993
timestamp 1663859327
transform 1 0 112560 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_111_996
timestamp 1663859327
transform 1 0 112896 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_111_1028
timestamp 1663859327
transform 1 0 116480 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_1044
timestamp 1663859327
transform 1 0 118272 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_2
timestamp 1663859327
transform 1 0 1568 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_112_7
timestamp 1663859327
transform 1 0 2128 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_112_23
timestamp 1663859327
transform 1 0 3920 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_31
timestamp 1663859327
transform 1 0 4816 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_37
timestamp 1663859327
transform 1 0 5488 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_101
timestamp 1663859327
transform 1 0 12656 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_105
timestamp 1663859327
transform 1 0 13104 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_108
timestamp 1663859327
transform 1 0 13440 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_172
timestamp 1663859327
transform 1 0 20608 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_176
timestamp 1663859327
transform 1 0 21056 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_179
timestamp 1663859327
transform 1 0 21392 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_243
timestamp 1663859327
transform 1 0 28560 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_247
timestamp 1663859327
transform 1 0 29008 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_250
timestamp 1663859327
transform 1 0 29344 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_314
timestamp 1663859327
transform 1 0 36512 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_318
timestamp 1663859327
transform 1 0 36960 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_321
timestamp 1663859327
transform 1 0 37296 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_385
timestamp 1663859327
transform 1 0 44464 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_389
timestamp 1663859327
transform 1 0 44912 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_392
timestamp 1663859327
transform 1 0 45248 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_456
timestamp 1663859327
transform 1 0 52416 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_460
timestamp 1663859327
transform 1 0 52864 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_463
timestamp 1663859327
transform 1 0 53200 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_527
timestamp 1663859327
transform 1 0 60368 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_531
timestamp 1663859327
transform 1 0 60816 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_534
timestamp 1663859327
transform 1 0 61152 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_598
timestamp 1663859327
transform 1 0 68320 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_602
timestamp 1663859327
transform 1 0 68768 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_605
timestamp 1663859327
transform 1 0 69104 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_669
timestamp 1663859327
transform 1 0 76272 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_673
timestamp 1663859327
transform 1 0 76720 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_676
timestamp 1663859327
transform 1 0 77056 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_740
timestamp 1663859327
transform 1 0 84224 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_744
timestamp 1663859327
transform 1 0 84672 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_747
timestamp 1663859327
transform 1 0 85008 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_811
timestamp 1663859327
transform 1 0 92176 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_815
timestamp 1663859327
transform 1 0 92624 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_818
timestamp 1663859327
transform 1 0 92960 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_882
timestamp 1663859327
transform 1 0 100128 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_886
timestamp 1663859327
transform 1 0 100576 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_889
timestamp 1663859327
transform 1 0 100912 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_953
timestamp 1663859327
transform 1 0 108080 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_957
timestamp 1663859327
transform 1 0 108528 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_960
timestamp 1663859327
transform 1 0 108864 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_1024
timestamp 1663859327
transform 1 0 116032 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1028
timestamp 1663859327
transform 1 0 116480 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_112_1031
timestamp 1663859327
transform 1 0 116816 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1039
timestamp 1663859327
transform 1 0 117712 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_1044
timestamp 1663859327
transform 1 0 118272 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_2
timestamp 1663859327
transform 1 0 1568 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_66
timestamp 1663859327
transform 1 0 8736 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_70
timestamp 1663859327
transform 1 0 9184 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_73
timestamp 1663859327
transform 1 0 9520 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_137
timestamp 1663859327
transform 1 0 16688 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_141
timestamp 1663859327
transform 1 0 17136 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_144
timestamp 1663859327
transform 1 0 17472 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_208
timestamp 1663859327
transform 1 0 24640 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_212
timestamp 1663859327
transform 1 0 25088 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_215
timestamp 1663859327
transform 1 0 25424 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_279
timestamp 1663859327
transform 1 0 32592 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_283
timestamp 1663859327
transform 1 0 33040 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_286
timestamp 1663859327
transform 1 0 33376 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_350
timestamp 1663859327
transform 1 0 40544 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_354
timestamp 1663859327
transform 1 0 40992 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_357
timestamp 1663859327
transform 1 0 41328 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_421
timestamp 1663859327
transform 1 0 48496 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_425
timestamp 1663859327
transform 1 0 48944 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_428
timestamp 1663859327
transform 1 0 49280 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_492
timestamp 1663859327
transform 1 0 56448 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_496
timestamp 1663859327
transform 1 0 56896 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_499
timestamp 1663859327
transform 1 0 57232 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_563
timestamp 1663859327
transform 1 0 64400 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_567
timestamp 1663859327
transform 1 0 64848 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_570
timestamp 1663859327
transform 1 0 65184 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_634
timestamp 1663859327
transform 1 0 72352 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_638
timestamp 1663859327
transform 1 0 72800 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_641
timestamp 1663859327
transform 1 0 73136 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_705
timestamp 1663859327
transform 1 0 80304 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_709
timestamp 1663859327
transform 1 0 80752 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_712
timestamp 1663859327
transform 1 0 81088 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_776
timestamp 1663859327
transform 1 0 88256 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_780
timestamp 1663859327
transform 1 0 88704 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_783
timestamp 1663859327
transform 1 0 89040 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_847
timestamp 1663859327
transform 1 0 96208 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_851
timestamp 1663859327
transform 1 0 96656 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_854
timestamp 1663859327
transform 1 0 96992 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_918
timestamp 1663859327
transform 1 0 104160 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_922
timestamp 1663859327
transform 1 0 104608 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_925
timestamp 1663859327
transform 1 0 104944 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_989
timestamp 1663859327
transform 1 0 112112 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_993
timestamp 1663859327
transform 1 0 112560 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_113_996
timestamp 1663859327
transform 1 0 112896 0 -1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_113_1028
timestamp 1663859327
transform 1 0 116480 0 -1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_1044
timestamp 1663859327
transform 1 0 118272 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_2
timestamp 1663859327
transform 1 0 1568 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_114_7
timestamp 1663859327
transform 1 0 2128 0 1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_114_23
timestamp 1663859327
transform 1 0 3920 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_31
timestamp 1663859327
transform 1 0 4816 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_37
timestamp 1663859327
transform 1 0 5488 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_101
timestamp 1663859327
transform 1 0 12656 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_105
timestamp 1663859327
transform 1 0 13104 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_108
timestamp 1663859327
transform 1 0 13440 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_172
timestamp 1663859327
transform 1 0 20608 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_176
timestamp 1663859327
transform 1 0 21056 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_179
timestamp 1663859327
transform 1 0 21392 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_243
timestamp 1663859327
transform 1 0 28560 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_247
timestamp 1663859327
transform 1 0 29008 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_250
timestamp 1663859327
transform 1 0 29344 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_314
timestamp 1663859327
transform 1 0 36512 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_318
timestamp 1663859327
transform 1 0 36960 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_321
timestamp 1663859327
transform 1 0 37296 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_385
timestamp 1663859327
transform 1 0 44464 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_389
timestamp 1663859327
transform 1 0 44912 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_392
timestamp 1663859327
transform 1 0 45248 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_456
timestamp 1663859327
transform 1 0 52416 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_460
timestamp 1663859327
transform 1 0 52864 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_463
timestamp 1663859327
transform 1 0 53200 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_527
timestamp 1663859327
transform 1 0 60368 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_531
timestamp 1663859327
transform 1 0 60816 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_534
timestamp 1663859327
transform 1 0 61152 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_598
timestamp 1663859327
transform 1 0 68320 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_602
timestamp 1663859327
transform 1 0 68768 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_605
timestamp 1663859327
transform 1 0 69104 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_669
timestamp 1663859327
transform 1 0 76272 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_673
timestamp 1663859327
transform 1 0 76720 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_676
timestamp 1663859327
transform 1 0 77056 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_740
timestamp 1663859327
transform 1 0 84224 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_744
timestamp 1663859327
transform 1 0 84672 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_747
timestamp 1663859327
transform 1 0 85008 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_811
timestamp 1663859327
transform 1 0 92176 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_815
timestamp 1663859327
transform 1 0 92624 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_818
timestamp 1663859327
transform 1 0 92960 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_882
timestamp 1663859327
transform 1 0 100128 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_886
timestamp 1663859327
transform 1 0 100576 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_889
timestamp 1663859327
transform 1 0 100912 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_953
timestamp 1663859327
transform 1 0 108080 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_957
timestamp 1663859327
transform 1 0 108528 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_960
timestamp 1663859327
transform 1 0 108864 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1024
timestamp 1663859327
transform 1 0 116032 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_1028
timestamp 1663859327
transform 1 0 116480 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_114_1031
timestamp 1663859327
transform 1 0 116816 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_1039
timestamp 1663859327
transform 1 0 117712 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_1043
timestamp 1663859327
transform 1 0 118160 0 1 92512
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_2
timestamp 1663859327
transform 1 0 1568 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_66
timestamp 1663859327
transform 1 0 8736 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_70
timestamp 1663859327
transform 1 0 9184 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_73
timestamp 1663859327
transform 1 0 9520 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_137
timestamp 1663859327
transform 1 0 16688 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_141
timestamp 1663859327
transform 1 0 17136 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_144
timestamp 1663859327
transform 1 0 17472 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_208
timestamp 1663859327
transform 1 0 24640 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_212
timestamp 1663859327
transform 1 0 25088 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_215
timestamp 1663859327
transform 1 0 25424 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_279
timestamp 1663859327
transform 1 0 32592 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_283
timestamp 1663859327
transform 1 0 33040 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_286
timestamp 1663859327
transform 1 0 33376 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_350
timestamp 1663859327
transform 1 0 40544 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_354
timestamp 1663859327
transform 1 0 40992 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_357
timestamp 1663859327
transform 1 0 41328 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_421
timestamp 1663859327
transform 1 0 48496 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_425
timestamp 1663859327
transform 1 0 48944 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_428
timestamp 1663859327
transform 1 0 49280 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_492
timestamp 1663859327
transform 1 0 56448 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_496
timestamp 1663859327
transform 1 0 56896 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_499
timestamp 1663859327
transform 1 0 57232 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_563
timestamp 1663859327
transform 1 0 64400 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_567
timestamp 1663859327
transform 1 0 64848 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_570
timestamp 1663859327
transform 1 0 65184 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_634
timestamp 1663859327
transform 1 0 72352 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_638
timestamp 1663859327
transform 1 0 72800 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_641
timestamp 1663859327
transform 1 0 73136 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_705
timestamp 1663859327
transform 1 0 80304 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_709
timestamp 1663859327
transform 1 0 80752 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_712
timestamp 1663859327
transform 1 0 81088 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_776
timestamp 1663859327
transform 1 0 88256 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_780
timestamp 1663859327
transform 1 0 88704 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_783
timestamp 1663859327
transform 1 0 89040 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_847
timestamp 1663859327
transform 1 0 96208 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_851
timestamp 1663859327
transform 1 0 96656 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_854
timestamp 1663859327
transform 1 0 96992 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_918
timestamp 1663859327
transform 1 0 104160 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_922
timestamp 1663859327
transform 1 0 104608 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_925
timestamp 1663859327
transform 1 0 104944 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_989
timestamp 1663859327
transform 1 0 112112 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_993
timestamp 1663859327
transform 1 0 112560 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_115_996
timestamp 1663859327
transform 1 0 112896 0 -1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_115_1028
timestamp 1663859327
transform 1 0 116480 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_1044
timestamp 1663859327
transform 1 0 118272 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_116_2
timestamp 1663859327
transform 1 0 1568 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_34
timestamp 1663859327
transform 1 0 5152 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_37
timestamp 1663859327
transform 1 0 5488 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_101
timestamp 1663859327
transform 1 0 12656 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_105
timestamp 1663859327
transform 1 0 13104 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_108
timestamp 1663859327
transform 1 0 13440 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_172
timestamp 1663859327
transform 1 0 20608 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_176
timestamp 1663859327
transform 1 0 21056 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_179
timestamp 1663859327
transform 1 0 21392 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_243
timestamp 1663859327
transform 1 0 28560 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_247
timestamp 1663859327
transform 1 0 29008 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_250
timestamp 1663859327
transform 1 0 29344 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_314
timestamp 1663859327
transform 1 0 36512 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_318
timestamp 1663859327
transform 1 0 36960 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_321
timestamp 1663859327
transform 1 0 37296 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_385
timestamp 1663859327
transform 1 0 44464 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_389
timestamp 1663859327
transform 1 0 44912 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_392
timestamp 1663859327
transform 1 0 45248 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_456
timestamp 1663859327
transform 1 0 52416 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_460
timestamp 1663859327
transform 1 0 52864 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_463
timestamp 1663859327
transform 1 0 53200 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_527
timestamp 1663859327
transform 1 0 60368 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_531
timestamp 1663859327
transform 1 0 60816 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_534
timestamp 1663859327
transform 1 0 61152 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_598
timestamp 1663859327
transform 1 0 68320 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_602
timestamp 1663859327
transform 1 0 68768 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_605
timestamp 1663859327
transform 1 0 69104 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_669
timestamp 1663859327
transform 1 0 76272 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_673
timestamp 1663859327
transform 1 0 76720 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_676
timestamp 1663859327
transform 1 0 77056 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_740
timestamp 1663859327
transform 1 0 84224 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_744
timestamp 1663859327
transform 1 0 84672 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_747
timestamp 1663859327
transform 1 0 85008 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_811
timestamp 1663859327
transform 1 0 92176 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_815
timestamp 1663859327
transform 1 0 92624 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_818
timestamp 1663859327
transform 1 0 92960 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_882
timestamp 1663859327
transform 1 0 100128 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_886
timestamp 1663859327
transform 1 0 100576 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_889
timestamp 1663859327
transform 1 0 100912 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_953
timestamp 1663859327
transform 1 0 108080 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_957
timestamp 1663859327
transform 1 0 108528 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_960
timestamp 1663859327
transform 1 0 108864 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1024
timestamp 1663859327
transform 1 0 116032 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_1028
timestamp 1663859327
transform 1 0 116480 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_116_1031
timestamp 1663859327
transform 1 0 116816 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_1039
timestamp 1663859327
transform 1 0 117712 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_116_1043
timestamp 1663859327
transform 1 0 118160 0 1 94080
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_2
timestamp 1663859327
transform 1 0 1568 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_7
timestamp 1663859327
transform 1 0 2128 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_73
timestamp 1663859327
transform 1 0 9520 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_137
timestamp 1663859327
transform 1 0 16688 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_141
timestamp 1663859327
transform 1 0 17136 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_144
timestamp 1663859327
transform 1 0 17472 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_208
timestamp 1663859327
transform 1 0 24640 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_212
timestamp 1663859327
transform 1 0 25088 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_215
timestamp 1663859327
transform 1 0 25424 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_279
timestamp 1663859327
transform 1 0 32592 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_283
timestamp 1663859327
transform 1 0 33040 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_286
timestamp 1663859327
transform 1 0 33376 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_350
timestamp 1663859327
transform 1 0 40544 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_354
timestamp 1663859327
transform 1 0 40992 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_357
timestamp 1663859327
transform 1 0 41328 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_421
timestamp 1663859327
transform 1 0 48496 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_425
timestamp 1663859327
transform 1 0 48944 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_428
timestamp 1663859327
transform 1 0 49280 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_492
timestamp 1663859327
transform 1 0 56448 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_496
timestamp 1663859327
transform 1 0 56896 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_499
timestamp 1663859327
transform 1 0 57232 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_563
timestamp 1663859327
transform 1 0 64400 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_567
timestamp 1663859327
transform 1 0 64848 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_570
timestamp 1663859327
transform 1 0 65184 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_634
timestamp 1663859327
transform 1 0 72352 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_638
timestamp 1663859327
transform 1 0 72800 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_641
timestamp 1663859327
transform 1 0 73136 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_705
timestamp 1663859327
transform 1 0 80304 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_709
timestamp 1663859327
transform 1 0 80752 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_712
timestamp 1663859327
transform 1 0 81088 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_776
timestamp 1663859327
transform 1 0 88256 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_780
timestamp 1663859327
transform 1 0 88704 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_783
timestamp 1663859327
transform 1 0 89040 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_847
timestamp 1663859327
transform 1 0 96208 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_851
timestamp 1663859327
transform 1 0 96656 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_854
timestamp 1663859327
transform 1 0 96992 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_918
timestamp 1663859327
transform 1 0 104160 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_922
timestamp 1663859327
transform 1 0 104608 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_925
timestamp 1663859327
transform 1 0 104944 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_989
timestamp 1663859327
transform 1 0 112112 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_993
timestamp 1663859327
transform 1 0 112560 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_117_996
timestamp 1663859327
transform 1 0 112896 0 -1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_117_1028
timestamp 1663859327
transform 1 0 116480 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_1044
timestamp 1663859327
transform 1 0 118272 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_2
timestamp 1663859327
transform 1 0 1568 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_34
timestamp 1663859327
transform 1 0 5152 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_37
timestamp 1663859327
transform 1 0 5488 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_101
timestamp 1663859327
transform 1 0 12656 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_105
timestamp 1663859327
transform 1 0 13104 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_108
timestamp 1663859327
transform 1 0 13440 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_172
timestamp 1663859327
transform 1 0 20608 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_176
timestamp 1663859327
transform 1 0 21056 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_179
timestamp 1663859327
transform 1 0 21392 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_243
timestamp 1663859327
transform 1 0 28560 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_247
timestamp 1663859327
transform 1 0 29008 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_250
timestamp 1663859327
transform 1 0 29344 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_314
timestamp 1663859327
transform 1 0 36512 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_318
timestamp 1663859327
transform 1 0 36960 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_321
timestamp 1663859327
transform 1 0 37296 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_385
timestamp 1663859327
transform 1 0 44464 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_389
timestamp 1663859327
transform 1 0 44912 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_392
timestamp 1663859327
transform 1 0 45248 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_456
timestamp 1663859327
transform 1 0 52416 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_460
timestamp 1663859327
transform 1 0 52864 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_463
timestamp 1663859327
transform 1 0 53200 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_527
timestamp 1663859327
transform 1 0 60368 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_531
timestamp 1663859327
transform 1 0 60816 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_534
timestamp 1663859327
transform 1 0 61152 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_598
timestamp 1663859327
transform 1 0 68320 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_602
timestamp 1663859327
transform 1 0 68768 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_605
timestamp 1663859327
transform 1 0 69104 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_669
timestamp 1663859327
transform 1 0 76272 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_673
timestamp 1663859327
transform 1 0 76720 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_676
timestamp 1663859327
transform 1 0 77056 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_740
timestamp 1663859327
transform 1 0 84224 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_744
timestamp 1663859327
transform 1 0 84672 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_747
timestamp 1663859327
transform 1 0 85008 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_811
timestamp 1663859327
transform 1 0 92176 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_815
timestamp 1663859327
transform 1 0 92624 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_818
timestamp 1663859327
transform 1 0 92960 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_882
timestamp 1663859327
transform 1 0 100128 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_886
timestamp 1663859327
transform 1 0 100576 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_889
timestamp 1663859327
transform 1 0 100912 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_953
timestamp 1663859327
transform 1 0 108080 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_957
timestamp 1663859327
transform 1 0 108528 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_118_960
timestamp 1663859327
transform 1 0 108864 0 1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_1024
timestamp 1663859327
transform 1 0 116032 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1028
timestamp 1663859327
transform 1 0 116480 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_1031
timestamp 1663859327
transform 1 0 116816 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1039
timestamp 1663859327
transform 1 0 117712 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_1044
timestamp 1663859327
transform 1 0 118272 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_2
timestamp 1663859327
transform 1 0 1568 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_7
timestamp 1663859327
transform 1 0 2128 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_73
timestamp 1663859327
transform 1 0 9520 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_137
timestamp 1663859327
transform 1 0 16688 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_141
timestamp 1663859327
transform 1 0 17136 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_144
timestamp 1663859327
transform 1 0 17472 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_208
timestamp 1663859327
transform 1 0 24640 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_212
timestamp 1663859327
transform 1 0 25088 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_215
timestamp 1663859327
transform 1 0 25424 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_279
timestamp 1663859327
transform 1 0 32592 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_283
timestamp 1663859327
transform 1 0 33040 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_286
timestamp 1663859327
transform 1 0 33376 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_350
timestamp 1663859327
transform 1 0 40544 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_354
timestamp 1663859327
transform 1 0 40992 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_357
timestamp 1663859327
transform 1 0 41328 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_421
timestamp 1663859327
transform 1 0 48496 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_425
timestamp 1663859327
transform 1 0 48944 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_428
timestamp 1663859327
transform 1 0 49280 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_492
timestamp 1663859327
transform 1 0 56448 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_496
timestamp 1663859327
transform 1 0 56896 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_499
timestamp 1663859327
transform 1 0 57232 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_563
timestamp 1663859327
transform 1 0 64400 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_567
timestamp 1663859327
transform 1 0 64848 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_570
timestamp 1663859327
transform 1 0 65184 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_634
timestamp 1663859327
transform 1 0 72352 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_638
timestamp 1663859327
transform 1 0 72800 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_641
timestamp 1663859327
transform 1 0 73136 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_705
timestamp 1663859327
transform 1 0 80304 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_709
timestamp 1663859327
transform 1 0 80752 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_712
timestamp 1663859327
transform 1 0 81088 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_776
timestamp 1663859327
transform 1 0 88256 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_780
timestamp 1663859327
transform 1 0 88704 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_783
timestamp 1663859327
transform 1 0 89040 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_847
timestamp 1663859327
transform 1 0 96208 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_851
timestamp 1663859327
transform 1 0 96656 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_854
timestamp 1663859327
transform 1 0 96992 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_918
timestamp 1663859327
transform 1 0 104160 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_922
timestamp 1663859327
transform 1 0 104608 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_119_925
timestamp 1663859327
transform 1 0 104944 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_989
timestamp 1663859327
transform 1 0 112112 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_993
timestamp 1663859327
transform 1 0 112560 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_119_996
timestamp 1663859327
transform 1 0 112896 0 -1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_119_1028
timestamp 1663859327
transform 1 0 116480 0 -1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_1044
timestamp 1663859327
transform 1 0 118272 0 -1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_120_2
timestamp 1663859327
transform 1 0 1568 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_34
timestamp 1663859327
transform 1 0 5152 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_37
timestamp 1663859327
transform 1 0 5488 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_101
timestamp 1663859327
transform 1 0 12656 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_105
timestamp 1663859327
transform 1 0 13104 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_108
timestamp 1663859327
transform 1 0 13440 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_172
timestamp 1663859327
transform 1 0 20608 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_176
timestamp 1663859327
transform 1 0 21056 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_179
timestamp 1663859327
transform 1 0 21392 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_243
timestamp 1663859327
transform 1 0 28560 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_247
timestamp 1663859327
transform 1 0 29008 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_250
timestamp 1663859327
transform 1 0 29344 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_314
timestamp 1663859327
transform 1 0 36512 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_318
timestamp 1663859327
transform 1 0 36960 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_321
timestamp 1663859327
transform 1 0 37296 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_385
timestamp 1663859327
transform 1 0 44464 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_389
timestamp 1663859327
transform 1 0 44912 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_392
timestamp 1663859327
transform 1 0 45248 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_456
timestamp 1663859327
transform 1 0 52416 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_460
timestamp 1663859327
transform 1 0 52864 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_463
timestamp 1663859327
transform 1 0 53200 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_527
timestamp 1663859327
transform 1 0 60368 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_531
timestamp 1663859327
transform 1 0 60816 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_534
timestamp 1663859327
transform 1 0 61152 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_598
timestamp 1663859327
transform 1 0 68320 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_602
timestamp 1663859327
transform 1 0 68768 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_605
timestamp 1663859327
transform 1 0 69104 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_669
timestamp 1663859327
transform 1 0 76272 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_673
timestamp 1663859327
transform 1 0 76720 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_676
timestamp 1663859327
transform 1 0 77056 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_740
timestamp 1663859327
transform 1 0 84224 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_744
timestamp 1663859327
transform 1 0 84672 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_747
timestamp 1663859327
transform 1 0 85008 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_811
timestamp 1663859327
transform 1 0 92176 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_815
timestamp 1663859327
transform 1 0 92624 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_818
timestamp 1663859327
transform 1 0 92960 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_882
timestamp 1663859327
transform 1 0 100128 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_886
timestamp 1663859327
transform 1 0 100576 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_889
timestamp 1663859327
transform 1 0 100912 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_953
timestamp 1663859327
transform 1 0 108080 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_957
timestamp 1663859327
transform 1 0 108528 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_120_960
timestamp 1663859327
transform 1 0 108864 0 1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_1024
timestamp 1663859327
transform 1 0 116032 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1028
timestamp 1663859327
transform 1 0 116480 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_120_1031
timestamp 1663859327
transform 1 0 116816 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1039
timestamp 1663859327
transform 1 0 117712 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_1044
timestamp 1663859327
transform 1 0 118272 0 1 97216
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_2
timestamp 1663859327
transform 1 0 1568 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_66
timestamp 1663859327
transform 1 0 8736 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_70
timestamp 1663859327
transform 1 0 9184 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_73
timestamp 1663859327
transform 1 0 9520 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_137
timestamp 1663859327
transform 1 0 16688 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_141
timestamp 1663859327
transform 1 0 17136 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_144
timestamp 1663859327
transform 1 0 17472 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_208
timestamp 1663859327
transform 1 0 24640 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_212
timestamp 1663859327
transform 1 0 25088 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_215
timestamp 1663859327
transform 1 0 25424 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_279
timestamp 1663859327
transform 1 0 32592 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_283
timestamp 1663859327
transform 1 0 33040 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_286
timestamp 1663859327
transform 1 0 33376 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_350
timestamp 1663859327
transform 1 0 40544 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_354
timestamp 1663859327
transform 1 0 40992 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_357
timestamp 1663859327
transform 1 0 41328 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_421
timestamp 1663859327
transform 1 0 48496 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_425
timestamp 1663859327
transform 1 0 48944 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_428
timestamp 1663859327
transform 1 0 49280 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_492
timestamp 1663859327
transform 1 0 56448 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_496
timestamp 1663859327
transform 1 0 56896 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_499
timestamp 1663859327
transform 1 0 57232 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_563
timestamp 1663859327
transform 1 0 64400 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_567
timestamp 1663859327
transform 1 0 64848 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_570
timestamp 1663859327
transform 1 0 65184 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_634
timestamp 1663859327
transform 1 0 72352 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_638
timestamp 1663859327
transform 1 0 72800 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_641
timestamp 1663859327
transform 1 0 73136 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_705
timestamp 1663859327
transform 1 0 80304 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_709
timestamp 1663859327
transform 1 0 80752 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_712
timestamp 1663859327
transform 1 0 81088 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_776
timestamp 1663859327
transform 1 0 88256 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_780
timestamp 1663859327
transform 1 0 88704 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_783
timestamp 1663859327
transform 1 0 89040 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_847
timestamp 1663859327
transform 1 0 96208 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_851
timestamp 1663859327
transform 1 0 96656 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_854
timestamp 1663859327
transform 1 0 96992 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_918
timestamp 1663859327
transform 1 0 104160 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_922
timestamp 1663859327
transform 1 0 104608 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_121_925
timestamp 1663859327
transform 1 0 104944 0 -1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_989
timestamp 1663859327
transform 1 0 112112 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_993
timestamp 1663859327
transform 1 0 112560 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_121_996
timestamp 1663859327
transform 1 0 112896 0 -1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_121_1028
timestamp 1663859327
transform 1 0 116480 0 -1 98784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_1036
timestamp 1663859327
transform 1 0 117376 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_1044
timestamp 1663859327
transform 1 0 118272 0 -1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_122_2
timestamp 1663859327
transform 1 0 1568 0 1 98784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_34
timestamp 1663859327
transform 1 0 5152 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_37
timestamp 1663859327
transform 1 0 5488 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_101
timestamp 1663859327
transform 1 0 12656 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_105
timestamp 1663859327
transform 1 0 13104 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_108
timestamp 1663859327
transform 1 0 13440 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_172
timestamp 1663859327
transform 1 0 20608 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_176
timestamp 1663859327
transform 1 0 21056 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_179
timestamp 1663859327
transform 1 0 21392 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_243
timestamp 1663859327
transform 1 0 28560 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_247
timestamp 1663859327
transform 1 0 29008 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_250
timestamp 1663859327
transform 1 0 29344 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_314
timestamp 1663859327
transform 1 0 36512 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_318
timestamp 1663859327
transform 1 0 36960 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_321
timestamp 1663859327
transform 1 0 37296 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_385
timestamp 1663859327
transform 1 0 44464 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_389
timestamp 1663859327
transform 1 0 44912 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_392
timestamp 1663859327
transform 1 0 45248 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_456
timestamp 1663859327
transform 1 0 52416 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_460
timestamp 1663859327
transform 1 0 52864 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_463
timestamp 1663859327
transform 1 0 53200 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_527
timestamp 1663859327
transform 1 0 60368 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_531
timestamp 1663859327
transform 1 0 60816 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_534
timestamp 1663859327
transform 1 0 61152 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_598
timestamp 1663859327
transform 1 0 68320 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_602
timestamp 1663859327
transform 1 0 68768 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_605
timestamp 1663859327
transform 1 0 69104 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_669
timestamp 1663859327
transform 1 0 76272 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_673
timestamp 1663859327
transform 1 0 76720 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_676
timestamp 1663859327
transform 1 0 77056 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_740
timestamp 1663859327
transform 1 0 84224 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_744
timestamp 1663859327
transform 1 0 84672 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_747
timestamp 1663859327
transform 1 0 85008 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_811
timestamp 1663859327
transform 1 0 92176 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_815
timestamp 1663859327
transform 1 0 92624 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_818
timestamp 1663859327
transform 1 0 92960 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_882
timestamp 1663859327
transform 1 0 100128 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_886
timestamp 1663859327
transform 1 0 100576 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_889
timestamp 1663859327
transform 1 0 100912 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_953
timestamp 1663859327
transform 1 0 108080 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_957
timestamp 1663859327
transform 1 0 108528 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_122_960
timestamp 1663859327
transform 1 0 108864 0 1 98784
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1024
timestamp 1663859327
transform 1 0 116032 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_1028
timestamp 1663859327
transform 1 0 116480 0 1 98784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_122_1031
timestamp 1663859327
transform 1 0 116816 0 1 98784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_1039
timestamp 1663859327
transform 1 0 117712 0 1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_122_1043
timestamp 1663859327
transform 1 0 118160 0 1 98784
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_2
timestamp 1663859327
transform 1 0 1568 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_66
timestamp 1663859327
transform 1 0 8736 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_70
timestamp 1663859327
transform 1 0 9184 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_73
timestamp 1663859327
transform 1 0 9520 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_137
timestamp 1663859327
transform 1 0 16688 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_141
timestamp 1663859327
transform 1 0 17136 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_144
timestamp 1663859327
transform 1 0 17472 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_208
timestamp 1663859327
transform 1 0 24640 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_212
timestamp 1663859327
transform 1 0 25088 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_215
timestamp 1663859327
transform 1 0 25424 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_279
timestamp 1663859327
transform 1 0 32592 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_283
timestamp 1663859327
transform 1 0 33040 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_286
timestamp 1663859327
transform 1 0 33376 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_350
timestamp 1663859327
transform 1 0 40544 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_354
timestamp 1663859327
transform 1 0 40992 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_357
timestamp 1663859327
transform 1 0 41328 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_421
timestamp 1663859327
transform 1 0 48496 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_425
timestamp 1663859327
transform 1 0 48944 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_428
timestamp 1663859327
transform 1 0 49280 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_492
timestamp 1663859327
transform 1 0 56448 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_496
timestamp 1663859327
transform 1 0 56896 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_499
timestamp 1663859327
transform 1 0 57232 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_563
timestamp 1663859327
transform 1 0 64400 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_567
timestamp 1663859327
transform 1 0 64848 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_570
timestamp 1663859327
transform 1 0 65184 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_634
timestamp 1663859327
transform 1 0 72352 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_638
timestamp 1663859327
transform 1 0 72800 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_641
timestamp 1663859327
transform 1 0 73136 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_705
timestamp 1663859327
transform 1 0 80304 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_709
timestamp 1663859327
transform 1 0 80752 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_712
timestamp 1663859327
transform 1 0 81088 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_776
timestamp 1663859327
transform 1 0 88256 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_780
timestamp 1663859327
transform 1 0 88704 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_783
timestamp 1663859327
transform 1 0 89040 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_847
timestamp 1663859327
transform 1 0 96208 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_851
timestamp 1663859327
transform 1 0 96656 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_854
timestamp 1663859327
transform 1 0 96992 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_918
timestamp 1663859327
transform 1 0 104160 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_922
timestamp 1663859327
transform 1 0 104608 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_123_925
timestamp 1663859327
transform 1 0 104944 0 -1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_989
timestamp 1663859327
transform 1 0 112112 0 -1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_993
timestamp 1663859327
transform 1 0 112560 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_123_996
timestamp 1663859327
transform 1 0 112896 0 -1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_123_1028
timestamp 1663859327
transform 1 0 116480 0 -1 100352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_1044
timestamp 1663859327
transform 1 0 118272 0 -1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_124_2
timestamp 1663859327
transform 1 0 1568 0 1 100352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_34
timestamp 1663859327
transform 1 0 5152 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_37
timestamp 1663859327
transform 1 0 5488 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_101
timestamp 1663859327
transform 1 0 12656 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_105
timestamp 1663859327
transform 1 0 13104 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_108
timestamp 1663859327
transform 1 0 13440 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_172
timestamp 1663859327
transform 1 0 20608 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_176
timestamp 1663859327
transform 1 0 21056 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_179
timestamp 1663859327
transform 1 0 21392 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_243
timestamp 1663859327
transform 1 0 28560 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_247
timestamp 1663859327
transform 1 0 29008 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_250
timestamp 1663859327
transform 1 0 29344 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_314
timestamp 1663859327
transform 1 0 36512 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_318
timestamp 1663859327
transform 1 0 36960 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_321
timestamp 1663859327
transform 1 0 37296 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_385
timestamp 1663859327
transform 1 0 44464 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_389
timestamp 1663859327
transform 1 0 44912 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_392
timestamp 1663859327
transform 1 0 45248 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_456
timestamp 1663859327
transform 1 0 52416 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_460
timestamp 1663859327
transform 1 0 52864 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_463
timestamp 1663859327
transform 1 0 53200 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_527
timestamp 1663859327
transform 1 0 60368 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_531
timestamp 1663859327
transform 1 0 60816 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_534
timestamp 1663859327
transform 1 0 61152 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_598
timestamp 1663859327
transform 1 0 68320 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_602
timestamp 1663859327
transform 1 0 68768 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_605
timestamp 1663859327
transform 1 0 69104 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_669
timestamp 1663859327
transform 1 0 76272 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_673
timestamp 1663859327
transform 1 0 76720 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_676
timestamp 1663859327
transform 1 0 77056 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_740
timestamp 1663859327
transform 1 0 84224 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_744
timestamp 1663859327
transform 1 0 84672 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_747
timestamp 1663859327
transform 1 0 85008 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_811
timestamp 1663859327
transform 1 0 92176 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_815
timestamp 1663859327
transform 1 0 92624 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_818
timestamp 1663859327
transform 1 0 92960 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_882
timestamp 1663859327
transform 1 0 100128 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_886
timestamp 1663859327
transform 1 0 100576 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_889
timestamp 1663859327
transform 1 0 100912 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_953
timestamp 1663859327
transform 1 0 108080 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_957
timestamp 1663859327
transform 1 0 108528 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_960
timestamp 1663859327
transform 1 0 108864 0 1 100352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1024
timestamp 1663859327
transform 1 0 116032 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_1028
timestamp 1663859327
transform 1 0 116480 0 1 100352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_124_1031
timestamp 1663859327
transform 1 0 116816 0 1 100352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_1039
timestamp 1663859327
transform 1 0 117712 0 1 100352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_124_1043
timestamp 1663859327
transform 1 0 118160 0 1 100352
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_2
timestamp 1663859327
transform 1 0 1568 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_7
timestamp 1663859327
transform 1 0 2128 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_73
timestamp 1663859327
transform 1 0 9520 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_137
timestamp 1663859327
transform 1 0 16688 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_141
timestamp 1663859327
transform 1 0 17136 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_144
timestamp 1663859327
transform 1 0 17472 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_208
timestamp 1663859327
transform 1 0 24640 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_212
timestamp 1663859327
transform 1 0 25088 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_215
timestamp 1663859327
transform 1 0 25424 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_279
timestamp 1663859327
transform 1 0 32592 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_283
timestamp 1663859327
transform 1 0 33040 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_286
timestamp 1663859327
transform 1 0 33376 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_350
timestamp 1663859327
transform 1 0 40544 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_354
timestamp 1663859327
transform 1 0 40992 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_357
timestamp 1663859327
transform 1 0 41328 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_421
timestamp 1663859327
transform 1 0 48496 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_425
timestamp 1663859327
transform 1 0 48944 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_428
timestamp 1663859327
transform 1 0 49280 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_492
timestamp 1663859327
transform 1 0 56448 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_496
timestamp 1663859327
transform 1 0 56896 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_499
timestamp 1663859327
transform 1 0 57232 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_563
timestamp 1663859327
transform 1 0 64400 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_567
timestamp 1663859327
transform 1 0 64848 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_570
timestamp 1663859327
transform 1 0 65184 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_634
timestamp 1663859327
transform 1 0 72352 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_638
timestamp 1663859327
transform 1 0 72800 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_641
timestamp 1663859327
transform 1 0 73136 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_705
timestamp 1663859327
transform 1 0 80304 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_709
timestamp 1663859327
transform 1 0 80752 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_712
timestamp 1663859327
transform 1 0 81088 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_776
timestamp 1663859327
transform 1 0 88256 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_780
timestamp 1663859327
transform 1 0 88704 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_783
timestamp 1663859327
transform 1 0 89040 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_847
timestamp 1663859327
transform 1 0 96208 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_851
timestamp 1663859327
transform 1 0 96656 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_854
timestamp 1663859327
transform 1 0 96992 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_918
timestamp 1663859327
transform 1 0 104160 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_922
timestamp 1663859327
transform 1 0 104608 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_125_925
timestamp 1663859327
transform 1 0 104944 0 -1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_989
timestamp 1663859327
transform 1 0 112112 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_993
timestamp 1663859327
transform 1 0 112560 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_125_996
timestamp 1663859327
transform 1 0 112896 0 -1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_125_1028
timestamp 1663859327
transform 1 0 116480 0 -1 101920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_1044
timestamp 1663859327
transform 1 0 118272 0 -1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_126_2
timestamp 1663859327
transform 1 0 1568 0 1 101920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_34
timestamp 1663859327
transform 1 0 5152 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_37
timestamp 1663859327
transform 1 0 5488 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_101
timestamp 1663859327
transform 1 0 12656 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_105
timestamp 1663859327
transform 1 0 13104 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_108
timestamp 1663859327
transform 1 0 13440 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_172
timestamp 1663859327
transform 1 0 20608 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_176
timestamp 1663859327
transform 1 0 21056 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_179
timestamp 1663859327
transform 1 0 21392 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_243
timestamp 1663859327
transform 1 0 28560 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_247
timestamp 1663859327
transform 1 0 29008 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_250
timestamp 1663859327
transform 1 0 29344 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_314
timestamp 1663859327
transform 1 0 36512 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_318
timestamp 1663859327
transform 1 0 36960 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_321
timestamp 1663859327
transform 1 0 37296 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_385
timestamp 1663859327
transform 1 0 44464 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_389
timestamp 1663859327
transform 1 0 44912 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_392
timestamp 1663859327
transform 1 0 45248 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_456
timestamp 1663859327
transform 1 0 52416 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_460
timestamp 1663859327
transform 1 0 52864 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_463
timestamp 1663859327
transform 1 0 53200 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_527
timestamp 1663859327
transform 1 0 60368 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_531
timestamp 1663859327
transform 1 0 60816 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_534
timestamp 1663859327
transform 1 0 61152 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_598
timestamp 1663859327
transform 1 0 68320 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_602
timestamp 1663859327
transform 1 0 68768 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_605
timestamp 1663859327
transform 1 0 69104 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_669
timestamp 1663859327
transform 1 0 76272 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_673
timestamp 1663859327
transform 1 0 76720 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_676
timestamp 1663859327
transform 1 0 77056 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_740
timestamp 1663859327
transform 1 0 84224 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_744
timestamp 1663859327
transform 1 0 84672 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_747
timestamp 1663859327
transform 1 0 85008 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_811
timestamp 1663859327
transform 1 0 92176 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_815
timestamp 1663859327
transform 1 0 92624 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_818
timestamp 1663859327
transform 1 0 92960 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_882
timestamp 1663859327
transform 1 0 100128 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_886
timestamp 1663859327
transform 1 0 100576 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_889
timestamp 1663859327
transform 1 0 100912 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_953
timestamp 1663859327
transform 1 0 108080 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_957
timestamp 1663859327
transform 1 0 108528 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_126_960
timestamp 1663859327
transform 1 0 108864 0 1 101920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1024
timestamp 1663859327
transform 1 0 116032 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_1028
timestamp 1663859327
transform 1 0 116480 0 1 101920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_126_1031
timestamp 1663859327
transform 1 0 116816 0 1 101920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_1039
timestamp 1663859327
transform 1 0 117712 0 1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_126_1043
timestamp 1663859327
transform 1 0 118160 0 1 101920
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_2
timestamp 1663859327
transform 1 0 1568 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_66
timestamp 1663859327
transform 1 0 8736 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_70
timestamp 1663859327
transform 1 0 9184 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_73
timestamp 1663859327
transform 1 0 9520 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_137
timestamp 1663859327
transform 1 0 16688 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_141
timestamp 1663859327
transform 1 0 17136 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_144
timestamp 1663859327
transform 1 0 17472 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_208
timestamp 1663859327
transform 1 0 24640 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_212
timestamp 1663859327
transform 1 0 25088 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_215
timestamp 1663859327
transform 1 0 25424 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_279
timestamp 1663859327
transform 1 0 32592 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_283
timestamp 1663859327
transform 1 0 33040 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_286
timestamp 1663859327
transform 1 0 33376 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_350
timestamp 1663859327
transform 1 0 40544 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_354
timestamp 1663859327
transform 1 0 40992 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_357
timestamp 1663859327
transform 1 0 41328 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_421
timestamp 1663859327
transform 1 0 48496 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_425
timestamp 1663859327
transform 1 0 48944 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_428
timestamp 1663859327
transform 1 0 49280 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_492
timestamp 1663859327
transform 1 0 56448 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_496
timestamp 1663859327
transform 1 0 56896 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_499
timestamp 1663859327
transform 1 0 57232 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_563
timestamp 1663859327
transform 1 0 64400 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_567
timestamp 1663859327
transform 1 0 64848 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_570
timestamp 1663859327
transform 1 0 65184 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_634
timestamp 1663859327
transform 1 0 72352 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_638
timestamp 1663859327
transform 1 0 72800 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_641
timestamp 1663859327
transform 1 0 73136 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_705
timestamp 1663859327
transform 1 0 80304 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_709
timestamp 1663859327
transform 1 0 80752 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_712
timestamp 1663859327
transform 1 0 81088 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_776
timestamp 1663859327
transform 1 0 88256 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_780
timestamp 1663859327
transform 1 0 88704 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_783
timestamp 1663859327
transform 1 0 89040 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_847
timestamp 1663859327
transform 1 0 96208 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_851
timestamp 1663859327
transform 1 0 96656 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_854
timestamp 1663859327
transform 1 0 96992 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_918
timestamp 1663859327
transform 1 0 104160 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_922
timestamp 1663859327
transform 1 0 104608 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_127_925
timestamp 1663859327
transform 1 0 104944 0 -1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_989
timestamp 1663859327
transform 1 0 112112 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_993
timestamp 1663859327
transform 1 0 112560 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_127_996
timestamp 1663859327
transform 1 0 112896 0 -1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_127_1028
timestamp 1663859327
transform 1 0 116480 0 -1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_1036
timestamp 1663859327
transform 1 0 117376 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_1044
timestamp 1663859327
transform 1 0 118272 0 -1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_128_2
timestamp 1663859327
transform 1 0 1568 0 1 103488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_34
timestamp 1663859327
transform 1 0 5152 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_37
timestamp 1663859327
transform 1 0 5488 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_101
timestamp 1663859327
transform 1 0 12656 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_105
timestamp 1663859327
transform 1 0 13104 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_108
timestamp 1663859327
transform 1 0 13440 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_172
timestamp 1663859327
transform 1 0 20608 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_176
timestamp 1663859327
transform 1 0 21056 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_179
timestamp 1663859327
transform 1 0 21392 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_243
timestamp 1663859327
transform 1 0 28560 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_247
timestamp 1663859327
transform 1 0 29008 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_250
timestamp 1663859327
transform 1 0 29344 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_314
timestamp 1663859327
transform 1 0 36512 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_318
timestamp 1663859327
transform 1 0 36960 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_321
timestamp 1663859327
transform 1 0 37296 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_385
timestamp 1663859327
transform 1 0 44464 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_389
timestamp 1663859327
transform 1 0 44912 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_392
timestamp 1663859327
transform 1 0 45248 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_456
timestamp 1663859327
transform 1 0 52416 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_460
timestamp 1663859327
transform 1 0 52864 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_463
timestamp 1663859327
transform 1 0 53200 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_527
timestamp 1663859327
transform 1 0 60368 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_531
timestamp 1663859327
transform 1 0 60816 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_534
timestamp 1663859327
transform 1 0 61152 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_598
timestamp 1663859327
transform 1 0 68320 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_602
timestamp 1663859327
transform 1 0 68768 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_605
timestamp 1663859327
transform 1 0 69104 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_669
timestamp 1663859327
transform 1 0 76272 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_673
timestamp 1663859327
transform 1 0 76720 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_676
timestamp 1663859327
transform 1 0 77056 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_740
timestamp 1663859327
transform 1 0 84224 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_744
timestamp 1663859327
transform 1 0 84672 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_747
timestamp 1663859327
transform 1 0 85008 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_811
timestamp 1663859327
transform 1 0 92176 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_815
timestamp 1663859327
transform 1 0 92624 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_818
timestamp 1663859327
transform 1 0 92960 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_882
timestamp 1663859327
transform 1 0 100128 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_886
timestamp 1663859327
transform 1 0 100576 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_889
timestamp 1663859327
transform 1 0 100912 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_953
timestamp 1663859327
transform 1 0 108080 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_957
timestamp 1663859327
transform 1 0 108528 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_960
timestamp 1663859327
transform 1 0 108864 0 1 103488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1024
timestamp 1663859327
transform 1 0 116032 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_1028
timestamp 1663859327
transform 1 0 116480 0 1 103488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_128_1031
timestamp 1663859327
transform 1 0 116816 0 1 103488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_1039
timestamp 1663859327
transform 1 0 117712 0 1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_128_1043
timestamp 1663859327
transform 1 0 118160 0 1 103488
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_2
timestamp 1663859327
transform 1 0 1568 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_66
timestamp 1663859327
transform 1 0 8736 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_70
timestamp 1663859327
transform 1 0 9184 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_73
timestamp 1663859327
transform 1 0 9520 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_137
timestamp 1663859327
transform 1 0 16688 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_141
timestamp 1663859327
transform 1 0 17136 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_144
timestamp 1663859327
transform 1 0 17472 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_208
timestamp 1663859327
transform 1 0 24640 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_212
timestamp 1663859327
transform 1 0 25088 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_215
timestamp 1663859327
transform 1 0 25424 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_279
timestamp 1663859327
transform 1 0 32592 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_283
timestamp 1663859327
transform 1 0 33040 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_286
timestamp 1663859327
transform 1 0 33376 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_350
timestamp 1663859327
transform 1 0 40544 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_354
timestamp 1663859327
transform 1 0 40992 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_357
timestamp 1663859327
transform 1 0 41328 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_421
timestamp 1663859327
transform 1 0 48496 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_425
timestamp 1663859327
transform 1 0 48944 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_428
timestamp 1663859327
transform 1 0 49280 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_492
timestamp 1663859327
transform 1 0 56448 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_496
timestamp 1663859327
transform 1 0 56896 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_499
timestamp 1663859327
transform 1 0 57232 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_563
timestamp 1663859327
transform 1 0 64400 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_567
timestamp 1663859327
transform 1 0 64848 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_570
timestamp 1663859327
transform 1 0 65184 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_634
timestamp 1663859327
transform 1 0 72352 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_638
timestamp 1663859327
transform 1 0 72800 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_641
timestamp 1663859327
transform 1 0 73136 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_705
timestamp 1663859327
transform 1 0 80304 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_709
timestamp 1663859327
transform 1 0 80752 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_712
timestamp 1663859327
transform 1 0 81088 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_776
timestamp 1663859327
transform 1 0 88256 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_780
timestamp 1663859327
transform 1 0 88704 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_783
timestamp 1663859327
transform 1 0 89040 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_847
timestamp 1663859327
transform 1 0 96208 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_851
timestamp 1663859327
transform 1 0 96656 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_854
timestamp 1663859327
transform 1 0 96992 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_918
timestamp 1663859327
transform 1 0 104160 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_922
timestamp 1663859327
transform 1 0 104608 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_129_925
timestamp 1663859327
transform 1 0 104944 0 -1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_989
timestamp 1663859327
transform 1 0 112112 0 -1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_993
timestamp 1663859327
transform 1 0 112560 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_129_996
timestamp 1663859327
transform 1 0 112896 0 -1 105056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_129_1028
timestamp 1663859327
transform 1 0 116480 0 -1 105056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_1044
timestamp 1663859327
transform 1 0 118272 0 -1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_2
timestamp 1663859327
transform 1 0 1568 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_130_7
timestamp 1663859327
transform 1 0 2128 0 1 105056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_130_23
timestamp 1663859327
transform 1 0 3920 0 1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_31
timestamp 1663859327
transform 1 0 4816 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_37
timestamp 1663859327
transform 1 0 5488 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_101
timestamp 1663859327
transform 1 0 12656 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_105
timestamp 1663859327
transform 1 0 13104 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_108
timestamp 1663859327
transform 1 0 13440 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_172
timestamp 1663859327
transform 1 0 20608 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_176
timestamp 1663859327
transform 1 0 21056 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_179
timestamp 1663859327
transform 1 0 21392 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_243
timestamp 1663859327
transform 1 0 28560 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_247
timestamp 1663859327
transform 1 0 29008 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_250
timestamp 1663859327
transform 1 0 29344 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_314
timestamp 1663859327
transform 1 0 36512 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_318
timestamp 1663859327
transform 1 0 36960 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_321
timestamp 1663859327
transform 1 0 37296 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_385
timestamp 1663859327
transform 1 0 44464 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_389
timestamp 1663859327
transform 1 0 44912 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_392
timestamp 1663859327
transform 1 0 45248 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_456
timestamp 1663859327
transform 1 0 52416 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_460
timestamp 1663859327
transform 1 0 52864 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_463
timestamp 1663859327
transform 1 0 53200 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_527
timestamp 1663859327
transform 1 0 60368 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_531
timestamp 1663859327
transform 1 0 60816 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_534
timestamp 1663859327
transform 1 0 61152 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_598
timestamp 1663859327
transform 1 0 68320 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_602
timestamp 1663859327
transform 1 0 68768 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_605
timestamp 1663859327
transform 1 0 69104 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_669
timestamp 1663859327
transform 1 0 76272 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_673
timestamp 1663859327
transform 1 0 76720 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_676
timestamp 1663859327
transform 1 0 77056 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_740
timestamp 1663859327
transform 1 0 84224 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_744
timestamp 1663859327
transform 1 0 84672 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_747
timestamp 1663859327
transform 1 0 85008 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_811
timestamp 1663859327
transform 1 0 92176 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_815
timestamp 1663859327
transform 1 0 92624 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_818
timestamp 1663859327
transform 1 0 92960 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_882
timestamp 1663859327
transform 1 0 100128 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_886
timestamp 1663859327
transform 1 0 100576 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_889
timestamp 1663859327
transform 1 0 100912 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_953
timestamp 1663859327
transform 1 0 108080 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_957
timestamp 1663859327
transform 1 0 108528 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_960
timestamp 1663859327
transform 1 0 108864 0 1 105056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1024
timestamp 1663859327
transform 1 0 116032 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_1028
timestamp 1663859327
transform 1 0 116480 0 1 105056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_130_1031
timestamp 1663859327
transform 1 0 116816 0 1 105056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_1039
timestamp 1663859327
transform 1 0 117712 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_130_1043
timestamp 1663859327
transform 1 0 118160 0 1 105056
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_2
timestamp 1663859327
transform 1 0 1568 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_66
timestamp 1663859327
transform 1 0 8736 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_70
timestamp 1663859327
transform 1 0 9184 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_73
timestamp 1663859327
transform 1 0 9520 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_137
timestamp 1663859327
transform 1 0 16688 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_141
timestamp 1663859327
transform 1 0 17136 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_144
timestamp 1663859327
transform 1 0 17472 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_208
timestamp 1663859327
transform 1 0 24640 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_212
timestamp 1663859327
transform 1 0 25088 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_215
timestamp 1663859327
transform 1 0 25424 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_279
timestamp 1663859327
transform 1 0 32592 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_283
timestamp 1663859327
transform 1 0 33040 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_286
timestamp 1663859327
transform 1 0 33376 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_350
timestamp 1663859327
transform 1 0 40544 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_354
timestamp 1663859327
transform 1 0 40992 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_357
timestamp 1663859327
transform 1 0 41328 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_421
timestamp 1663859327
transform 1 0 48496 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_425
timestamp 1663859327
transform 1 0 48944 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_428
timestamp 1663859327
transform 1 0 49280 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_492
timestamp 1663859327
transform 1 0 56448 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_496
timestamp 1663859327
transform 1 0 56896 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_499
timestamp 1663859327
transform 1 0 57232 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_563
timestamp 1663859327
transform 1 0 64400 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_567
timestamp 1663859327
transform 1 0 64848 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_570
timestamp 1663859327
transform 1 0 65184 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_634
timestamp 1663859327
transform 1 0 72352 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_638
timestamp 1663859327
transform 1 0 72800 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_641
timestamp 1663859327
transform 1 0 73136 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_705
timestamp 1663859327
transform 1 0 80304 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_709
timestamp 1663859327
transform 1 0 80752 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_712
timestamp 1663859327
transform 1 0 81088 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_776
timestamp 1663859327
transform 1 0 88256 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_780
timestamp 1663859327
transform 1 0 88704 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_783
timestamp 1663859327
transform 1 0 89040 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_847
timestamp 1663859327
transform 1 0 96208 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_851
timestamp 1663859327
transform 1 0 96656 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_854
timestamp 1663859327
transform 1 0 96992 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_918
timestamp 1663859327
transform 1 0 104160 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_922
timestamp 1663859327
transform 1 0 104608 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_131_925
timestamp 1663859327
transform 1 0 104944 0 -1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_989
timestamp 1663859327
transform 1 0 112112 0 -1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_993
timestamp 1663859327
transform 1 0 112560 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_131_996
timestamp 1663859327
transform 1 0 112896 0 -1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_131_1028
timestamp 1663859327
transform 1 0 116480 0 -1 106624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_1044
timestamp 1663859327
transform 1 0 118272 0 -1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_132_2
timestamp 1663859327
transform 1 0 1568 0 1 106624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_34
timestamp 1663859327
transform 1 0 5152 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_37
timestamp 1663859327
transform 1 0 5488 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_101
timestamp 1663859327
transform 1 0 12656 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_105
timestamp 1663859327
transform 1 0 13104 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_108
timestamp 1663859327
transform 1 0 13440 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_172
timestamp 1663859327
transform 1 0 20608 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_176
timestamp 1663859327
transform 1 0 21056 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_179
timestamp 1663859327
transform 1 0 21392 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_243
timestamp 1663859327
transform 1 0 28560 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_247
timestamp 1663859327
transform 1 0 29008 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_250
timestamp 1663859327
transform 1 0 29344 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_314
timestamp 1663859327
transform 1 0 36512 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_318
timestamp 1663859327
transform 1 0 36960 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_321
timestamp 1663859327
transform 1 0 37296 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_385
timestamp 1663859327
transform 1 0 44464 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_389
timestamp 1663859327
transform 1 0 44912 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_392
timestamp 1663859327
transform 1 0 45248 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_456
timestamp 1663859327
transform 1 0 52416 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_460
timestamp 1663859327
transform 1 0 52864 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_463
timestamp 1663859327
transform 1 0 53200 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_527
timestamp 1663859327
transform 1 0 60368 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_531
timestamp 1663859327
transform 1 0 60816 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_534
timestamp 1663859327
transform 1 0 61152 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_598
timestamp 1663859327
transform 1 0 68320 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_602
timestamp 1663859327
transform 1 0 68768 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_605
timestamp 1663859327
transform 1 0 69104 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_669
timestamp 1663859327
transform 1 0 76272 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_673
timestamp 1663859327
transform 1 0 76720 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_676
timestamp 1663859327
transform 1 0 77056 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_740
timestamp 1663859327
transform 1 0 84224 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_744
timestamp 1663859327
transform 1 0 84672 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_747
timestamp 1663859327
transform 1 0 85008 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_811
timestamp 1663859327
transform 1 0 92176 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_815
timestamp 1663859327
transform 1 0 92624 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_818
timestamp 1663859327
transform 1 0 92960 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_882
timestamp 1663859327
transform 1 0 100128 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_886
timestamp 1663859327
transform 1 0 100576 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_889
timestamp 1663859327
transform 1 0 100912 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_953
timestamp 1663859327
transform 1 0 108080 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_957
timestamp 1663859327
transform 1 0 108528 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_960
timestamp 1663859327
transform 1 0 108864 0 1 106624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_1024
timestamp 1663859327
transform 1 0 116032 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1028
timestamp 1663859327
transform 1 0 116480 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_132_1031
timestamp 1663859327
transform 1 0 116816 0 1 106624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1039
timestamp 1663859327
transform 1 0 117712 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_1044
timestamp 1663859327
transform 1 0 118272 0 1 106624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_2
timestamp 1663859327
transform 1 0 1568 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_66
timestamp 1663859327
transform 1 0 8736 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_70
timestamp 1663859327
transform 1 0 9184 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_73
timestamp 1663859327
transform 1 0 9520 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_137
timestamp 1663859327
transform 1 0 16688 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_141
timestamp 1663859327
transform 1 0 17136 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_144
timestamp 1663859327
transform 1 0 17472 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_208
timestamp 1663859327
transform 1 0 24640 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_212
timestamp 1663859327
transform 1 0 25088 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_215
timestamp 1663859327
transform 1 0 25424 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_279
timestamp 1663859327
transform 1 0 32592 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_283
timestamp 1663859327
transform 1 0 33040 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_286
timestamp 1663859327
transform 1 0 33376 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_350
timestamp 1663859327
transform 1 0 40544 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_354
timestamp 1663859327
transform 1 0 40992 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_357
timestamp 1663859327
transform 1 0 41328 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_421
timestamp 1663859327
transform 1 0 48496 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_425
timestamp 1663859327
transform 1 0 48944 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_428
timestamp 1663859327
transform 1 0 49280 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_492
timestamp 1663859327
transform 1 0 56448 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_496
timestamp 1663859327
transform 1 0 56896 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_499
timestamp 1663859327
transform 1 0 57232 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_563
timestamp 1663859327
transform 1 0 64400 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_567
timestamp 1663859327
transform 1 0 64848 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_570
timestamp 1663859327
transform 1 0 65184 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_634
timestamp 1663859327
transform 1 0 72352 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_638
timestamp 1663859327
transform 1 0 72800 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_641
timestamp 1663859327
transform 1 0 73136 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_705
timestamp 1663859327
transform 1 0 80304 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_709
timestamp 1663859327
transform 1 0 80752 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_712
timestamp 1663859327
transform 1 0 81088 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_776
timestamp 1663859327
transform 1 0 88256 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_780
timestamp 1663859327
transform 1 0 88704 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_783
timestamp 1663859327
transform 1 0 89040 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_847
timestamp 1663859327
transform 1 0 96208 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_851
timestamp 1663859327
transform 1 0 96656 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_854
timestamp 1663859327
transform 1 0 96992 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_918
timestamp 1663859327
transform 1 0 104160 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_922
timestamp 1663859327
transform 1 0 104608 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_133_925
timestamp 1663859327
transform 1 0 104944 0 -1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_989
timestamp 1663859327
transform 1 0 112112 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_993
timestamp 1663859327
transform 1 0 112560 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_133_996
timestamp 1663859327
transform 1 0 112896 0 -1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_133_1028
timestamp 1663859327
transform 1 0 116480 0 -1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_1036
timestamp 1663859327
transform 1 0 117376 0 -1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_1044
timestamp 1663859327
transform 1 0 118272 0 -1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_134_2
timestamp 1663859327
transform 1 0 1568 0 1 108192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_34
timestamp 1663859327
transform 1 0 5152 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_37
timestamp 1663859327
transform 1 0 5488 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_101
timestamp 1663859327
transform 1 0 12656 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_105
timestamp 1663859327
transform 1 0 13104 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_108
timestamp 1663859327
transform 1 0 13440 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_172
timestamp 1663859327
transform 1 0 20608 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_176
timestamp 1663859327
transform 1 0 21056 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_179
timestamp 1663859327
transform 1 0 21392 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_243
timestamp 1663859327
transform 1 0 28560 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_247
timestamp 1663859327
transform 1 0 29008 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_250
timestamp 1663859327
transform 1 0 29344 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_314
timestamp 1663859327
transform 1 0 36512 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_318
timestamp 1663859327
transform 1 0 36960 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_321
timestamp 1663859327
transform 1 0 37296 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_385
timestamp 1663859327
transform 1 0 44464 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_389
timestamp 1663859327
transform 1 0 44912 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_392
timestamp 1663859327
transform 1 0 45248 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_456
timestamp 1663859327
transform 1 0 52416 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_460
timestamp 1663859327
transform 1 0 52864 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_463
timestamp 1663859327
transform 1 0 53200 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_527
timestamp 1663859327
transform 1 0 60368 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_531
timestamp 1663859327
transform 1 0 60816 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_534
timestamp 1663859327
transform 1 0 61152 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_598
timestamp 1663859327
transform 1 0 68320 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_602
timestamp 1663859327
transform 1 0 68768 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_605
timestamp 1663859327
transform 1 0 69104 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_669
timestamp 1663859327
transform 1 0 76272 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_673
timestamp 1663859327
transform 1 0 76720 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_676
timestamp 1663859327
transform 1 0 77056 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_740
timestamp 1663859327
transform 1 0 84224 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_744
timestamp 1663859327
transform 1 0 84672 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_747
timestamp 1663859327
transform 1 0 85008 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_811
timestamp 1663859327
transform 1 0 92176 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_815
timestamp 1663859327
transform 1 0 92624 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_818
timestamp 1663859327
transform 1 0 92960 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_882
timestamp 1663859327
transform 1 0 100128 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_886
timestamp 1663859327
transform 1 0 100576 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_889
timestamp 1663859327
transform 1 0 100912 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_953
timestamp 1663859327
transform 1 0 108080 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_957
timestamp 1663859327
transform 1 0 108528 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_960
timestamp 1663859327
transform 1 0 108864 0 1 108192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1024
timestamp 1663859327
transform 1 0 116032 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_1028
timestamp 1663859327
transform 1 0 116480 0 1 108192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_134_1031
timestamp 1663859327
transform 1 0 116816 0 1 108192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_1039
timestamp 1663859327
transform 1 0 117712 0 1 108192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_134_1043
timestamp 1663859327
transform 1 0 118160 0 1 108192
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_2
timestamp 1663859327
transform 1 0 1568 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_66
timestamp 1663859327
transform 1 0 8736 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_70
timestamp 1663859327
transform 1 0 9184 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_73
timestamp 1663859327
transform 1 0 9520 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_137
timestamp 1663859327
transform 1 0 16688 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_141
timestamp 1663859327
transform 1 0 17136 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_144
timestamp 1663859327
transform 1 0 17472 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_208
timestamp 1663859327
transform 1 0 24640 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_212
timestamp 1663859327
transform 1 0 25088 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_215
timestamp 1663859327
transform 1 0 25424 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_279
timestamp 1663859327
transform 1 0 32592 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_283
timestamp 1663859327
transform 1 0 33040 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_286
timestamp 1663859327
transform 1 0 33376 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_350
timestamp 1663859327
transform 1 0 40544 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_354
timestamp 1663859327
transform 1 0 40992 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_357
timestamp 1663859327
transform 1 0 41328 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_421
timestamp 1663859327
transform 1 0 48496 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_425
timestamp 1663859327
transform 1 0 48944 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_428
timestamp 1663859327
transform 1 0 49280 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_492
timestamp 1663859327
transform 1 0 56448 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_496
timestamp 1663859327
transform 1 0 56896 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_499
timestamp 1663859327
transform 1 0 57232 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_563
timestamp 1663859327
transform 1 0 64400 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_567
timestamp 1663859327
transform 1 0 64848 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_570
timestamp 1663859327
transform 1 0 65184 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_634
timestamp 1663859327
transform 1 0 72352 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_638
timestamp 1663859327
transform 1 0 72800 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_641
timestamp 1663859327
transform 1 0 73136 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_705
timestamp 1663859327
transform 1 0 80304 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_709
timestamp 1663859327
transform 1 0 80752 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_712
timestamp 1663859327
transform 1 0 81088 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_776
timestamp 1663859327
transform 1 0 88256 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_780
timestamp 1663859327
transform 1 0 88704 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_783
timestamp 1663859327
transform 1 0 89040 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_847
timestamp 1663859327
transform 1 0 96208 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_851
timestamp 1663859327
transform 1 0 96656 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_854
timestamp 1663859327
transform 1 0 96992 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_918
timestamp 1663859327
transform 1 0 104160 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_922
timestamp 1663859327
transform 1 0 104608 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_135_925
timestamp 1663859327
transform 1 0 104944 0 -1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_989
timestamp 1663859327
transform 1 0 112112 0 -1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_993
timestamp 1663859327
transform 1 0 112560 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_135_996
timestamp 1663859327
transform 1 0 112896 0 -1 109760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_135_1028
timestamp 1663859327
transform 1 0 116480 0 -1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_1044
timestamp 1663859327
transform 1 0 118272 0 -1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_2
timestamp 1663859327
transform 1 0 1568 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_136_7
timestamp 1663859327
transform 1 0 2128 0 1 109760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_136_23
timestamp 1663859327
transform 1 0 3920 0 1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_31
timestamp 1663859327
transform 1 0 4816 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_37
timestamp 1663859327
transform 1 0 5488 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_101
timestamp 1663859327
transform 1 0 12656 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_105
timestamp 1663859327
transform 1 0 13104 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_108
timestamp 1663859327
transform 1 0 13440 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_172
timestamp 1663859327
transform 1 0 20608 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_176
timestamp 1663859327
transform 1 0 21056 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_179
timestamp 1663859327
transform 1 0 21392 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_243
timestamp 1663859327
transform 1 0 28560 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_247
timestamp 1663859327
transform 1 0 29008 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_250
timestamp 1663859327
transform 1 0 29344 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_314
timestamp 1663859327
transform 1 0 36512 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_318
timestamp 1663859327
transform 1 0 36960 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_321
timestamp 1663859327
transform 1 0 37296 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_385
timestamp 1663859327
transform 1 0 44464 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_389
timestamp 1663859327
transform 1 0 44912 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_392
timestamp 1663859327
transform 1 0 45248 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_456
timestamp 1663859327
transform 1 0 52416 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_460
timestamp 1663859327
transform 1 0 52864 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_463
timestamp 1663859327
transform 1 0 53200 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_527
timestamp 1663859327
transform 1 0 60368 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_531
timestamp 1663859327
transform 1 0 60816 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_534
timestamp 1663859327
transform 1 0 61152 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_598
timestamp 1663859327
transform 1 0 68320 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_602
timestamp 1663859327
transform 1 0 68768 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_605
timestamp 1663859327
transform 1 0 69104 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_669
timestamp 1663859327
transform 1 0 76272 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_673
timestamp 1663859327
transform 1 0 76720 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_676
timestamp 1663859327
transform 1 0 77056 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_740
timestamp 1663859327
transform 1 0 84224 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_744
timestamp 1663859327
transform 1 0 84672 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_747
timestamp 1663859327
transform 1 0 85008 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_811
timestamp 1663859327
transform 1 0 92176 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_815
timestamp 1663859327
transform 1 0 92624 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_818
timestamp 1663859327
transform 1 0 92960 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_882
timestamp 1663859327
transform 1 0 100128 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_886
timestamp 1663859327
transform 1 0 100576 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_889
timestamp 1663859327
transform 1 0 100912 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_953
timestamp 1663859327
transform 1 0 108080 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_957
timestamp 1663859327
transform 1 0 108528 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_136_960
timestamp 1663859327
transform 1 0 108864 0 1 109760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1024
timestamp 1663859327
transform 1 0 116032 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_1028
timestamp 1663859327
transform 1 0 116480 0 1 109760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_136_1031
timestamp 1663859327
transform 1 0 116816 0 1 109760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_1039
timestamp 1663859327
transform 1 0 117712 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_136_1043
timestamp 1663859327
transform 1 0 118160 0 1 109760
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_2
timestamp 1663859327
transform 1 0 1568 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_66
timestamp 1663859327
transform 1 0 8736 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_70
timestamp 1663859327
transform 1 0 9184 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_73
timestamp 1663859327
transform 1 0 9520 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_137
timestamp 1663859327
transform 1 0 16688 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_141
timestamp 1663859327
transform 1 0 17136 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_144
timestamp 1663859327
transform 1 0 17472 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_208
timestamp 1663859327
transform 1 0 24640 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_212
timestamp 1663859327
transform 1 0 25088 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_215
timestamp 1663859327
transform 1 0 25424 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_279
timestamp 1663859327
transform 1 0 32592 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_283
timestamp 1663859327
transform 1 0 33040 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_286
timestamp 1663859327
transform 1 0 33376 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_350
timestamp 1663859327
transform 1 0 40544 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_354
timestamp 1663859327
transform 1 0 40992 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_357
timestamp 1663859327
transform 1 0 41328 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_421
timestamp 1663859327
transform 1 0 48496 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_425
timestamp 1663859327
transform 1 0 48944 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_428
timestamp 1663859327
transform 1 0 49280 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_492
timestamp 1663859327
transform 1 0 56448 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_496
timestamp 1663859327
transform 1 0 56896 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_499
timestamp 1663859327
transform 1 0 57232 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_563
timestamp 1663859327
transform 1 0 64400 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_567
timestamp 1663859327
transform 1 0 64848 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_570
timestamp 1663859327
transform 1 0 65184 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_634
timestamp 1663859327
transform 1 0 72352 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_638
timestamp 1663859327
transform 1 0 72800 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_641
timestamp 1663859327
transform 1 0 73136 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_705
timestamp 1663859327
transform 1 0 80304 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_709
timestamp 1663859327
transform 1 0 80752 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_712
timestamp 1663859327
transform 1 0 81088 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_776
timestamp 1663859327
transform 1 0 88256 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_780
timestamp 1663859327
transform 1 0 88704 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_783
timestamp 1663859327
transform 1 0 89040 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_847
timestamp 1663859327
transform 1 0 96208 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_851
timestamp 1663859327
transform 1 0 96656 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_854
timestamp 1663859327
transform 1 0 96992 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_918
timestamp 1663859327
transform 1 0 104160 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_922
timestamp 1663859327
transform 1 0 104608 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_137_925
timestamp 1663859327
transform 1 0 104944 0 -1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_989
timestamp 1663859327
transform 1 0 112112 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_993
timestamp 1663859327
transform 1 0 112560 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_137_996
timestamp 1663859327
transform 1 0 112896 0 -1 111328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_137_1028
timestamp 1663859327
transform 1 0 116480 0 -1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_1036
timestamp 1663859327
transform 1 0 117376 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_1044
timestamp 1663859327
transform 1 0 118272 0 -1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_2
timestamp 1663859327
transform 1 0 1568 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_138_7
timestamp 1663859327
transform 1 0 2128 0 1 111328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_138_23
timestamp 1663859327
transform 1 0 3920 0 1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_31
timestamp 1663859327
transform 1 0 4816 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_37
timestamp 1663859327
transform 1 0 5488 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_101
timestamp 1663859327
transform 1 0 12656 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_105
timestamp 1663859327
transform 1 0 13104 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_108
timestamp 1663859327
transform 1 0 13440 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_172
timestamp 1663859327
transform 1 0 20608 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_176
timestamp 1663859327
transform 1 0 21056 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_179
timestamp 1663859327
transform 1 0 21392 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_243
timestamp 1663859327
transform 1 0 28560 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_247
timestamp 1663859327
transform 1 0 29008 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_250
timestamp 1663859327
transform 1 0 29344 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_314
timestamp 1663859327
transform 1 0 36512 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_318
timestamp 1663859327
transform 1 0 36960 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_321
timestamp 1663859327
transform 1 0 37296 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_385
timestamp 1663859327
transform 1 0 44464 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_389
timestamp 1663859327
transform 1 0 44912 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_392
timestamp 1663859327
transform 1 0 45248 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_456
timestamp 1663859327
transform 1 0 52416 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_460
timestamp 1663859327
transform 1 0 52864 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_463
timestamp 1663859327
transform 1 0 53200 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_527
timestamp 1663859327
transform 1 0 60368 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_531
timestamp 1663859327
transform 1 0 60816 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_534
timestamp 1663859327
transform 1 0 61152 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_598
timestamp 1663859327
transform 1 0 68320 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_602
timestamp 1663859327
transform 1 0 68768 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_605
timestamp 1663859327
transform 1 0 69104 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_669
timestamp 1663859327
transform 1 0 76272 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_673
timestamp 1663859327
transform 1 0 76720 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_676
timestamp 1663859327
transform 1 0 77056 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_740
timestamp 1663859327
transform 1 0 84224 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_744
timestamp 1663859327
transform 1 0 84672 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_747
timestamp 1663859327
transform 1 0 85008 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_811
timestamp 1663859327
transform 1 0 92176 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_815
timestamp 1663859327
transform 1 0 92624 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_818
timestamp 1663859327
transform 1 0 92960 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_882
timestamp 1663859327
transform 1 0 100128 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_886
timestamp 1663859327
transform 1 0 100576 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_889
timestamp 1663859327
transform 1 0 100912 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_953
timestamp 1663859327
transform 1 0 108080 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_957
timestamp 1663859327
transform 1 0 108528 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_138_960
timestamp 1663859327
transform 1 0 108864 0 1 111328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_1024
timestamp 1663859327
transform 1 0 116032 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1028
timestamp 1663859327
transform 1 0 116480 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_138_1031
timestamp 1663859327
transform 1 0 116816 0 1 111328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1039
timestamp 1663859327
transform 1 0 117712 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_1044
timestamp 1663859327
transform 1 0 118272 0 1 111328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_2
timestamp 1663859327
transform 1 0 1568 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_66
timestamp 1663859327
transform 1 0 8736 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_70
timestamp 1663859327
transform 1 0 9184 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_73
timestamp 1663859327
transform 1 0 9520 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_137
timestamp 1663859327
transform 1 0 16688 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_141
timestamp 1663859327
transform 1 0 17136 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_144
timestamp 1663859327
transform 1 0 17472 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_208
timestamp 1663859327
transform 1 0 24640 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_212
timestamp 1663859327
transform 1 0 25088 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_215
timestamp 1663859327
transform 1 0 25424 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_279
timestamp 1663859327
transform 1 0 32592 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_283
timestamp 1663859327
transform 1 0 33040 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_286
timestamp 1663859327
transform 1 0 33376 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_350
timestamp 1663859327
transform 1 0 40544 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_354
timestamp 1663859327
transform 1 0 40992 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_357
timestamp 1663859327
transform 1 0 41328 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_421
timestamp 1663859327
transform 1 0 48496 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_425
timestamp 1663859327
transform 1 0 48944 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_428
timestamp 1663859327
transform 1 0 49280 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_492
timestamp 1663859327
transform 1 0 56448 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_496
timestamp 1663859327
transform 1 0 56896 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_499
timestamp 1663859327
transform 1 0 57232 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_563
timestamp 1663859327
transform 1 0 64400 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_567
timestamp 1663859327
transform 1 0 64848 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_570
timestamp 1663859327
transform 1 0 65184 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_634
timestamp 1663859327
transform 1 0 72352 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_638
timestamp 1663859327
transform 1 0 72800 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_641
timestamp 1663859327
transform 1 0 73136 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_705
timestamp 1663859327
transform 1 0 80304 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_709
timestamp 1663859327
transform 1 0 80752 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_712
timestamp 1663859327
transform 1 0 81088 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_776
timestamp 1663859327
transform 1 0 88256 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_780
timestamp 1663859327
transform 1 0 88704 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_783
timestamp 1663859327
transform 1 0 89040 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_847
timestamp 1663859327
transform 1 0 96208 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_851
timestamp 1663859327
transform 1 0 96656 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_854
timestamp 1663859327
transform 1 0 96992 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_918
timestamp 1663859327
transform 1 0 104160 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_922
timestamp 1663859327
transform 1 0 104608 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_139_925
timestamp 1663859327
transform 1 0 104944 0 -1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_989
timestamp 1663859327
transform 1 0 112112 0 -1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_993
timestamp 1663859327
transform 1 0 112560 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_139_996
timestamp 1663859327
transform 1 0 112896 0 -1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_139_1028
timestamp 1663859327
transform 1 0 116480 0 -1 112896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_1044
timestamp 1663859327
transform 1 0 118272 0 -1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_140_2
timestamp 1663859327
transform 1 0 1568 0 1 112896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_34
timestamp 1663859327
transform 1 0 5152 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_37
timestamp 1663859327
transform 1 0 5488 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_101
timestamp 1663859327
transform 1 0 12656 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_105
timestamp 1663859327
transform 1 0 13104 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_108
timestamp 1663859327
transform 1 0 13440 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_172
timestamp 1663859327
transform 1 0 20608 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_176
timestamp 1663859327
transform 1 0 21056 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_179
timestamp 1663859327
transform 1 0 21392 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_243
timestamp 1663859327
transform 1 0 28560 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_247
timestamp 1663859327
transform 1 0 29008 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_250
timestamp 1663859327
transform 1 0 29344 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_314
timestamp 1663859327
transform 1 0 36512 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_318
timestamp 1663859327
transform 1 0 36960 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_321
timestamp 1663859327
transform 1 0 37296 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_385
timestamp 1663859327
transform 1 0 44464 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_389
timestamp 1663859327
transform 1 0 44912 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_392
timestamp 1663859327
transform 1 0 45248 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_456
timestamp 1663859327
transform 1 0 52416 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_460
timestamp 1663859327
transform 1 0 52864 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_463
timestamp 1663859327
transform 1 0 53200 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_527
timestamp 1663859327
transform 1 0 60368 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_531
timestamp 1663859327
transform 1 0 60816 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_534
timestamp 1663859327
transform 1 0 61152 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_598
timestamp 1663859327
transform 1 0 68320 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_602
timestamp 1663859327
transform 1 0 68768 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_605
timestamp 1663859327
transform 1 0 69104 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_669
timestamp 1663859327
transform 1 0 76272 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_673
timestamp 1663859327
transform 1 0 76720 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_676
timestamp 1663859327
transform 1 0 77056 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_740
timestamp 1663859327
transform 1 0 84224 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_744
timestamp 1663859327
transform 1 0 84672 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_747
timestamp 1663859327
transform 1 0 85008 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_811
timestamp 1663859327
transform 1 0 92176 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_815
timestamp 1663859327
transform 1 0 92624 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_818
timestamp 1663859327
transform 1 0 92960 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_882
timestamp 1663859327
transform 1 0 100128 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_886
timestamp 1663859327
transform 1 0 100576 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_889
timestamp 1663859327
transform 1 0 100912 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_953
timestamp 1663859327
transform 1 0 108080 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_957
timestamp 1663859327
transform 1 0 108528 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_140_960
timestamp 1663859327
transform 1 0 108864 0 1 112896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1024
timestamp 1663859327
transform 1 0 116032 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_1028
timestamp 1663859327
transform 1 0 116480 0 1 112896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_140_1031
timestamp 1663859327
transform 1 0 116816 0 1 112896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_1039
timestamp 1663859327
transform 1 0 117712 0 1 112896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_140_1043
timestamp 1663859327
transform 1 0 118160 0 1 112896
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_2
timestamp 1663859327
transform 1 0 1568 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_66
timestamp 1663859327
transform 1 0 8736 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_70
timestamp 1663859327
transform 1 0 9184 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_73
timestamp 1663859327
transform 1 0 9520 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_137
timestamp 1663859327
transform 1 0 16688 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_141
timestamp 1663859327
transform 1 0 17136 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_144
timestamp 1663859327
transform 1 0 17472 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_208
timestamp 1663859327
transform 1 0 24640 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_212
timestamp 1663859327
transform 1 0 25088 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_215
timestamp 1663859327
transform 1 0 25424 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_279
timestamp 1663859327
transform 1 0 32592 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_283
timestamp 1663859327
transform 1 0 33040 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_286
timestamp 1663859327
transform 1 0 33376 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_350
timestamp 1663859327
transform 1 0 40544 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_354
timestamp 1663859327
transform 1 0 40992 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_357
timestamp 1663859327
transform 1 0 41328 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_421
timestamp 1663859327
transform 1 0 48496 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_425
timestamp 1663859327
transform 1 0 48944 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_428
timestamp 1663859327
transform 1 0 49280 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_492
timestamp 1663859327
transform 1 0 56448 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_496
timestamp 1663859327
transform 1 0 56896 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_499
timestamp 1663859327
transform 1 0 57232 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_563
timestamp 1663859327
transform 1 0 64400 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_567
timestamp 1663859327
transform 1 0 64848 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_570
timestamp 1663859327
transform 1 0 65184 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_634
timestamp 1663859327
transform 1 0 72352 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_638
timestamp 1663859327
transform 1 0 72800 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_641
timestamp 1663859327
transform 1 0 73136 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_705
timestamp 1663859327
transform 1 0 80304 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_709
timestamp 1663859327
transform 1 0 80752 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_712
timestamp 1663859327
transform 1 0 81088 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_776
timestamp 1663859327
transform 1 0 88256 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_780
timestamp 1663859327
transform 1 0 88704 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_783
timestamp 1663859327
transform 1 0 89040 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_847
timestamp 1663859327
transform 1 0 96208 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_851
timestamp 1663859327
transform 1 0 96656 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_854
timestamp 1663859327
transform 1 0 96992 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_918
timestamp 1663859327
transform 1 0 104160 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_922
timestamp 1663859327
transform 1 0 104608 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_141_925
timestamp 1663859327
transform 1 0 104944 0 -1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_989
timestamp 1663859327
transform 1 0 112112 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_993
timestamp 1663859327
transform 1 0 112560 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_141_996
timestamp 1663859327
transform 1 0 112896 0 -1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_141_1028
timestamp 1663859327
transform 1 0 116480 0 -1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_141_1036
timestamp 1663859327
transform 1 0 117376 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_1044
timestamp 1663859327
transform 1 0 118272 0 -1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_142_2
timestamp 1663859327
transform 1 0 1568 0 1 114464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_34
timestamp 1663859327
transform 1 0 5152 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_37
timestamp 1663859327
transform 1 0 5488 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_101
timestamp 1663859327
transform 1 0 12656 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_105
timestamp 1663859327
transform 1 0 13104 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_108
timestamp 1663859327
transform 1 0 13440 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_172
timestamp 1663859327
transform 1 0 20608 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_176
timestamp 1663859327
transform 1 0 21056 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_179
timestamp 1663859327
transform 1 0 21392 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_243
timestamp 1663859327
transform 1 0 28560 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_247
timestamp 1663859327
transform 1 0 29008 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_250
timestamp 1663859327
transform 1 0 29344 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_314
timestamp 1663859327
transform 1 0 36512 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_318
timestamp 1663859327
transform 1 0 36960 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_321
timestamp 1663859327
transform 1 0 37296 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_385
timestamp 1663859327
transform 1 0 44464 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_389
timestamp 1663859327
transform 1 0 44912 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_392
timestamp 1663859327
transform 1 0 45248 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_456
timestamp 1663859327
transform 1 0 52416 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_460
timestamp 1663859327
transform 1 0 52864 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_463
timestamp 1663859327
transform 1 0 53200 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_527
timestamp 1663859327
transform 1 0 60368 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_531
timestamp 1663859327
transform 1 0 60816 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_534
timestamp 1663859327
transform 1 0 61152 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_598
timestamp 1663859327
transform 1 0 68320 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_602
timestamp 1663859327
transform 1 0 68768 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_605
timestamp 1663859327
transform 1 0 69104 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_669
timestamp 1663859327
transform 1 0 76272 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_673
timestamp 1663859327
transform 1 0 76720 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_676
timestamp 1663859327
transform 1 0 77056 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_740
timestamp 1663859327
transform 1 0 84224 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_744
timestamp 1663859327
transform 1 0 84672 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_747
timestamp 1663859327
transform 1 0 85008 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_811
timestamp 1663859327
transform 1 0 92176 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_815
timestamp 1663859327
transform 1 0 92624 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_818
timestamp 1663859327
transform 1 0 92960 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_882
timestamp 1663859327
transform 1 0 100128 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_886
timestamp 1663859327
transform 1 0 100576 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_889
timestamp 1663859327
transform 1 0 100912 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_953
timestamp 1663859327
transform 1 0 108080 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_957
timestamp 1663859327
transform 1 0 108528 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_142_960
timestamp 1663859327
transform 1 0 108864 0 1 114464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1024
timestamp 1663859327
transform 1 0 116032 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_1028
timestamp 1663859327
transform 1 0 116480 0 1 114464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_142_1031
timestamp 1663859327
transform 1 0 116816 0 1 114464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_1039
timestamp 1663859327
transform 1 0 117712 0 1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_1043
timestamp 1663859327
transform 1 0 118160 0 1 114464
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_2
timestamp 1663859327
transform 1 0 1568 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_66
timestamp 1663859327
transform 1 0 8736 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_70
timestamp 1663859327
transform 1 0 9184 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_73
timestamp 1663859327
transform 1 0 9520 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_137
timestamp 1663859327
transform 1 0 16688 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_141
timestamp 1663859327
transform 1 0 17136 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_144
timestamp 1663859327
transform 1 0 17472 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_208
timestamp 1663859327
transform 1 0 24640 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_212
timestamp 1663859327
transform 1 0 25088 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_215
timestamp 1663859327
transform 1 0 25424 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_279
timestamp 1663859327
transform 1 0 32592 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_283
timestamp 1663859327
transform 1 0 33040 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_286
timestamp 1663859327
transform 1 0 33376 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_350
timestamp 1663859327
transform 1 0 40544 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_354
timestamp 1663859327
transform 1 0 40992 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_357
timestamp 1663859327
transform 1 0 41328 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_421
timestamp 1663859327
transform 1 0 48496 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_425
timestamp 1663859327
transform 1 0 48944 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_428
timestamp 1663859327
transform 1 0 49280 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_492
timestamp 1663859327
transform 1 0 56448 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_496
timestamp 1663859327
transform 1 0 56896 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_499
timestamp 1663859327
transform 1 0 57232 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_563
timestamp 1663859327
transform 1 0 64400 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_567
timestamp 1663859327
transform 1 0 64848 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_570
timestamp 1663859327
transform 1 0 65184 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_634
timestamp 1663859327
transform 1 0 72352 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_638
timestamp 1663859327
transform 1 0 72800 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_641
timestamp 1663859327
transform 1 0 73136 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_705
timestamp 1663859327
transform 1 0 80304 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_709
timestamp 1663859327
transform 1 0 80752 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_712
timestamp 1663859327
transform 1 0 81088 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_776
timestamp 1663859327
transform 1 0 88256 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_780
timestamp 1663859327
transform 1 0 88704 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_783
timestamp 1663859327
transform 1 0 89040 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_847
timestamp 1663859327
transform 1 0 96208 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_851
timestamp 1663859327
transform 1 0 96656 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_854
timestamp 1663859327
transform 1 0 96992 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_918
timestamp 1663859327
transform 1 0 104160 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_922
timestamp 1663859327
transform 1 0 104608 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_143_925
timestamp 1663859327
transform 1 0 104944 0 -1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_989
timestamp 1663859327
transform 1 0 112112 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_993
timestamp 1663859327
transform 1 0 112560 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_143_996
timestamp 1663859327
transform 1 0 112896 0 -1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_143_1028
timestamp 1663859327
transform 1 0 116480 0 -1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_1036
timestamp 1663859327
transform 1 0 117376 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_1044
timestamp 1663859327
transform 1 0 118272 0 -1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_144_2
timestamp 1663859327
transform 1 0 1568 0 1 116032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_34
timestamp 1663859327
transform 1 0 5152 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_37
timestamp 1663859327
transform 1 0 5488 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_101
timestamp 1663859327
transform 1 0 12656 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_105
timestamp 1663859327
transform 1 0 13104 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_108
timestamp 1663859327
transform 1 0 13440 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_172
timestamp 1663859327
transform 1 0 20608 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_176
timestamp 1663859327
transform 1 0 21056 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_179
timestamp 1663859327
transform 1 0 21392 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_243
timestamp 1663859327
transform 1 0 28560 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_247
timestamp 1663859327
transform 1 0 29008 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_250
timestamp 1663859327
transform 1 0 29344 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_314
timestamp 1663859327
transform 1 0 36512 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_318
timestamp 1663859327
transform 1 0 36960 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_321
timestamp 1663859327
transform 1 0 37296 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_385
timestamp 1663859327
transform 1 0 44464 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_389
timestamp 1663859327
transform 1 0 44912 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_392
timestamp 1663859327
transform 1 0 45248 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_456
timestamp 1663859327
transform 1 0 52416 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_460
timestamp 1663859327
transform 1 0 52864 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_463
timestamp 1663859327
transform 1 0 53200 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_527
timestamp 1663859327
transform 1 0 60368 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_531
timestamp 1663859327
transform 1 0 60816 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_534
timestamp 1663859327
transform 1 0 61152 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_598
timestamp 1663859327
transform 1 0 68320 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_602
timestamp 1663859327
transform 1 0 68768 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_605
timestamp 1663859327
transform 1 0 69104 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_669
timestamp 1663859327
transform 1 0 76272 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_673
timestamp 1663859327
transform 1 0 76720 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_676
timestamp 1663859327
transform 1 0 77056 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_740
timestamp 1663859327
transform 1 0 84224 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_744
timestamp 1663859327
transform 1 0 84672 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_747
timestamp 1663859327
transform 1 0 85008 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_811
timestamp 1663859327
transform 1 0 92176 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_815
timestamp 1663859327
transform 1 0 92624 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_818
timestamp 1663859327
transform 1 0 92960 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_882
timestamp 1663859327
transform 1 0 100128 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_886
timestamp 1663859327
transform 1 0 100576 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_889
timestamp 1663859327
transform 1 0 100912 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_953
timestamp 1663859327
transform 1 0 108080 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_957
timestamp 1663859327
transform 1 0 108528 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_144_960
timestamp 1663859327
transform 1 0 108864 0 1 116032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_144_1024
timestamp 1663859327
transform 1 0 116032 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1028
timestamp 1663859327
transform 1 0 116480 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_144_1031
timestamp 1663859327
transform 1 0 116816 0 1 116032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1039
timestamp 1663859327
transform 1 0 117712 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_144_1044
timestamp 1663859327
transform 1 0 118272 0 1 116032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_2
timestamp 1663859327
transform 1 0 1568 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_7
timestamp 1663859327
transform 1 0 2128 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_73
timestamp 1663859327
transform 1 0 9520 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_137
timestamp 1663859327
transform 1 0 16688 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_141
timestamp 1663859327
transform 1 0 17136 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_144
timestamp 1663859327
transform 1 0 17472 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_208
timestamp 1663859327
transform 1 0 24640 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_212
timestamp 1663859327
transform 1 0 25088 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_215
timestamp 1663859327
transform 1 0 25424 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_279
timestamp 1663859327
transform 1 0 32592 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_283
timestamp 1663859327
transform 1 0 33040 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_286
timestamp 1663859327
transform 1 0 33376 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_350
timestamp 1663859327
transform 1 0 40544 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_354
timestamp 1663859327
transform 1 0 40992 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_357
timestamp 1663859327
transform 1 0 41328 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_421
timestamp 1663859327
transform 1 0 48496 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_425
timestamp 1663859327
transform 1 0 48944 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_428
timestamp 1663859327
transform 1 0 49280 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_492
timestamp 1663859327
transform 1 0 56448 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_496
timestamp 1663859327
transform 1 0 56896 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_499
timestamp 1663859327
transform 1 0 57232 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_563
timestamp 1663859327
transform 1 0 64400 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_567
timestamp 1663859327
transform 1 0 64848 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_570
timestamp 1663859327
transform 1 0 65184 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_634
timestamp 1663859327
transform 1 0 72352 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_638
timestamp 1663859327
transform 1 0 72800 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_641
timestamp 1663859327
transform 1 0 73136 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_705
timestamp 1663859327
transform 1 0 80304 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_709
timestamp 1663859327
transform 1 0 80752 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_712
timestamp 1663859327
transform 1 0 81088 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_776
timestamp 1663859327
transform 1 0 88256 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_780
timestamp 1663859327
transform 1 0 88704 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_783
timestamp 1663859327
transform 1 0 89040 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_847
timestamp 1663859327
transform 1 0 96208 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_851
timestamp 1663859327
transform 1 0 96656 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_854
timestamp 1663859327
transform 1 0 96992 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_918
timestamp 1663859327
transform 1 0 104160 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_922
timestamp 1663859327
transform 1 0 104608 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_145_925
timestamp 1663859327
transform 1 0 104944 0 -1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_145_989
timestamp 1663859327
transform 1 0 112112 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_993
timestamp 1663859327
transform 1 0 112560 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_145_996
timestamp 1663859327
transform 1 0 112896 0 -1 117600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_145_1028
timestamp 1663859327
transform 1 0 116480 0 -1 117600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_145_1044
timestamp 1663859327
transform 1 0 118272 0 -1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_146_2
timestamp 1663859327
transform 1 0 1568 0 1 117600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_34
timestamp 1663859327
transform 1 0 5152 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_37
timestamp 1663859327
transform 1 0 5488 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_101
timestamp 1663859327
transform 1 0 12656 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_105
timestamp 1663859327
transform 1 0 13104 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_108
timestamp 1663859327
transform 1 0 13440 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_172
timestamp 1663859327
transform 1 0 20608 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_176
timestamp 1663859327
transform 1 0 21056 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_179
timestamp 1663859327
transform 1 0 21392 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_243
timestamp 1663859327
transform 1 0 28560 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_247
timestamp 1663859327
transform 1 0 29008 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_250
timestamp 1663859327
transform 1 0 29344 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_314
timestamp 1663859327
transform 1 0 36512 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_318
timestamp 1663859327
transform 1 0 36960 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_321
timestamp 1663859327
transform 1 0 37296 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_385
timestamp 1663859327
transform 1 0 44464 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_389
timestamp 1663859327
transform 1 0 44912 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_392
timestamp 1663859327
transform 1 0 45248 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_456
timestamp 1663859327
transform 1 0 52416 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_460
timestamp 1663859327
transform 1 0 52864 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_463
timestamp 1663859327
transform 1 0 53200 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_527
timestamp 1663859327
transform 1 0 60368 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_531
timestamp 1663859327
transform 1 0 60816 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_534
timestamp 1663859327
transform 1 0 61152 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_598
timestamp 1663859327
transform 1 0 68320 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_602
timestamp 1663859327
transform 1 0 68768 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_605
timestamp 1663859327
transform 1 0 69104 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_669
timestamp 1663859327
transform 1 0 76272 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_673
timestamp 1663859327
transform 1 0 76720 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_676
timestamp 1663859327
transform 1 0 77056 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_740
timestamp 1663859327
transform 1 0 84224 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_744
timestamp 1663859327
transform 1 0 84672 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_747
timestamp 1663859327
transform 1 0 85008 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_811
timestamp 1663859327
transform 1 0 92176 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_815
timestamp 1663859327
transform 1 0 92624 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_818
timestamp 1663859327
transform 1 0 92960 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_882
timestamp 1663859327
transform 1 0 100128 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_886
timestamp 1663859327
transform 1 0 100576 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_889
timestamp 1663859327
transform 1 0 100912 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_953
timestamp 1663859327
transform 1 0 108080 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_957
timestamp 1663859327
transform 1 0 108528 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_146_960
timestamp 1663859327
transform 1 0 108864 0 1 117600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_1024
timestamp 1663859327
transform 1 0 116032 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_146_1028
timestamp 1663859327
transform 1 0 116480 0 1 117600
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_146_1031
timestamp 1663859327
transform 1 0 116816 0 1 117600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_146_1039
timestamp 1663859327
transform 1 0 117712 0 1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_146_1043
timestamp 1663859327
transform 1 0 118160 0 1 117600
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_2
timestamp 1663859327
transform 1 0 1568 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_66
timestamp 1663859327
transform 1 0 8736 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_70
timestamp 1663859327
transform 1 0 9184 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_73
timestamp 1663859327
transform 1 0 9520 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_137
timestamp 1663859327
transform 1 0 16688 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_141
timestamp 1663859327
transform 1 0 17136 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_144
timestamp 1663859327
transform 1 0 17472 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_208
timestamp 1663859327
transform 1 0 24640 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_212
timestamp 1663859327
transform 1 0 25088 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_215
timestamp 1663859327
transform 1 0 25424 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_279
timestamp 1663859327
transform 1 0 32592 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_283
timestamp 1663859327
transform 1 0 33040 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_286
timestamp 1663859327
transform 1 0 33376 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_350
timestamp 1663859327
transform 1 0 40544 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_354
timestamp 1663859327
transform 1 0 40992 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_357
timestamp 1663859327
transform 1 0 41328 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_421
timestamp 1663859327
transform 1 0 48496 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_425
timestamp 1663859327
transform 1 0 48944 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_428
timestamp 1663859327
transform 1 0 49280 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_492
timestamp 1663859327
transform 1 0 56448 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_496
timestamp 1663859327
transform 1 0 56896 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_499
timestamp 1663859327
transform 1 0 57232 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_563
timestamp 1663859327
transform 1 0 64400 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_567
timestamp 1663859327
transform 1 0 64848 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_570
timestamp 1663859327
transform 1 0 65184 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_634
timestamp 1663859327
transform 1 0 72352 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_638
timestamp 1663859327
transform 1 0 72800 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_641
timestamp 1663859327
transform 1 0 73136 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_705
timestamp 1663859327
transform 1 0 80304 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_709
timestamp 1663859327
transform 1 0 80752 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_712
timestamp 1663859327
transform 1 0 81088 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_776
timestamp 1663859327
transform 1 0 88256 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_780
timestamp 1663859327
transform 1 0 88704 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_783
timestamp 1663859327
transform 1 0 89040 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_847
timestamp 1663859327
transform 1 0 96208 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_851
timestamp 1663859327
transform 1 0 96656 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_854
timestamp 1663859327
transform 1 0 96992 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_918
timestamp 1663859327
transform 1 0 104160 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_922
timestamp 1663859327
transform 1 0 104608 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_147_925
timestamp 1663859327
transform 1 0 104944 0 -1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_147_989
timestamp 1663859327
transform 1 0 112112 0 -1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_993
timestamp 1663859327
transform 1 0 112560 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_147_996
timestamp 1663859327
transform 1 0 112896 0 -1 119168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_147_1028
timestamp 1663859327
transform 1 0 116480 0 -1 119168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_147_1044
timestamp 1663859327
transform 1 0 118272 0 -1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_148_2
timestamp 1663859327
transform 1 0 1568 0 1 119168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_34
timestamp 1663859327
transform 1 0 5152 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_37
timestamp 1663859327
transform 1 0 5488 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_101
timestamp 1663859327
transform 1 0 12656 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_105
timestamp 1663859327
transform 1 0 13104 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_108
timestamp 1663859327
transform 1 0 13440 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_172
timestamp 1663859327
transform 1 0 20608 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_176
timestamp 1663859327
transform 1 0 21056 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_179
timestamp 1663859327
transform 1 0 21392 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_243
timestamp 1663859327
transform 1 0 28560 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_247
timestamp 1663859327
transform 1 0 29008 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_250
timestamp 1663859327
transform 1 0 29344 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_314
timestamp 1663859327
transform 1 0 36512 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_318
timestamp 1663859327
transform 1 0 36960 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_321
timestamp 1663859327
transform 1 0 37296 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_385
timestamp 1663859327
transform 1 0 44464 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_389
timestamp 1663859327
transform 1 0 44912 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_392
timestamp 1663859327
transform 1 0 45248 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_456
timestamp 1663859327
transform 1 0 52416 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_460
timestamp 1663859327
transform 1 0 52864 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_463
timestamp 1663859327
transform 1 0 53200 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_527
timestamp 1663859327
transform 1 0 60368 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_531
timestamp 1663859327
transform 1 0 60816 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_534
timestamp 1663859327
transform 1 0 61152 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_598
timestamp 1663859327
transform 1 0 68320 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_602
timestamp 1663859327
transform 1 0 68768 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_605
timestamp 1663859327
transform 1 0 69104 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_669
timestamp 1663859327
transform 1 0 76272 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_673
timestamp 1663859327
transform 1 0 76720 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_676
timestamp 1663859327
transform 1 0 77056 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_740
timestamp 1663859327
transform 1 0 84224 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_744
timestamp 1663859327
transform 1 0 84672 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_747
timestamp 1663859327
transform 1 0 85008 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_811
timestamp 1663859327
transform 1 0 92176 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_815
timestamp 1663859327
transform 1 0 92624 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_818
timestamp 1663859327
transform 1 0 92960 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_882
timestamp 1663859327
transform 1 0 100128 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_886
timestamp 1663859327
transform 1 0 100576 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_889
timestamp 1663859327
transform 1 0 100912 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_953
timestamp 1663859327
transform 1 0 108080 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_957
timestamp 1663859327
transform 1 0 108528 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_148_960
timestamp 1663859327
transform 1 0 108864 0 1 119168
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_1024
timestamp 1663859327
transform 1 0 116032 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_148_1028
timestamp 1663859327
transform 1 0 116480 0 1 119168
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_148_1031
timestamp 1663859327
transform 1 0 116816 0 1 119168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_148_1039
timestamp 1663859327
transform 1 0 117712 0 1 119168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_148_1043
timestamp 1663859327
transform 1 0 118160 0 1 119168
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_2
timestamp 1663859327
transform 1 0 1568 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_66
timestamp 1663859327
transform 1 0 8736 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_70
timestamp 1663859327
transform 1 0 9184 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_73
timestamp 1663859327
transform 1 0 9520 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_137
timestamp 1663859327
transform 1 0 16688 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_141
timestamp 1663859327
transform 1 0 17136 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_144
timestamp 1663859327
transform 1 0 17472 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_208
timestamp 1663859327
transform 1 0 24640 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_212
timestamp 1663859327
transform 1 0 25088 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_215
timestamp 1663859327
transform 1 0 25424 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_279
timestamp 1663859327
transform 1 0 32592 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_283
timestamp 1663859327
transform 1 0 33040 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_286
timestamp 1663859327
transform 1 0 33376 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_350
timestamp 1663859327
transform 1 0 40544 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_354
timestamp 1663859327
transform 1 0 40992 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_357
timestamp 1663859327
transform 1 0 41328 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_421
timestamp 1663859327
transform 1 0 48496 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_425
timestamp 1663859327
transform 1 0 48944 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_428
timestamp 1663859327
transform 1 0 49280 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_492
timestamp 1663859327
transform 1 0 56448 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_496
timestamp 1663859327
transform 1 0 56896 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_499
timestamp 1663859327
transform 1 0 57232 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_563
timestamp 1663859327
transform 1 0 64400 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_567
timestamp 1663859327
transform 1 0 64848 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_570
timestamp 1663859327
transform 1 0 65184 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_634
timestamp 1663859327
transform 1 0 72352 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_638
timestamp 1663859327
transform 1 0 72800 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_641
timestamp 1663859327
transform 1 0 73136 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_705
timestamp 1663859327
transform 1 0 80304 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_709
timestamp 1663859327
transform 1 0 80752 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_712
timestamp 1663859327
transform 1 0 81088 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_776
timestamp 1663859327
transform 1 0 88256 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_780
timestamp 1663859327
transform 1 0 88704 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_783
timestamp 1663859327
transform 1 0 89040 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_847
timestamp 1663859327
transform 1 0 96208 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_851
timestamp 1663859327
transform 1 0 96656 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_854
timestamp 1663859327
transform 1 0 96992 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_918
timestamp 1663859327
transform 1 0 104160 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_922
timestamp 1663859327
transform 1 0 104608 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_149_925
timestamp 1663859327
transform 1 0 104944 0 -1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_149_989
timestamp 1663859327
transform 1 0 112112 0 -1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_993
timestamp 1663859327
transform 1 0 112560 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_149_996
timestamp 1663859327
transform 1 0 112896 0 -1 120736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_149_1028
timestamp 1663859327
transform 1 0 116480 0 -1 120736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_149_1044
timestamp 1663859327
transform 1 0 118272 0 -1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_150_2
timestamp 1663859327
transform 1 0 1568 0 1 120736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_34
timestamp 1663859327
transform 1 0 5152 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_37
timestamp 1663859327
transform 1 0 5488 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_101
timestamp 1663859327
transform 1 0 12656 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_105
timestamp 1663859327
transform 1 0 13104 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_108
timestamp 1663859327
transform 1 0 13440 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_172
timestamp 1663859327
transform 1 0 20608 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_176
timestamp 1663859327
transform 1 0 21056 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_179
timestamp 1663859327
transform 1 0 21392 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_243
timestamp 1663859327
transform 1 0 28560 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_247
timestamp 1663859327
transform 1 0 29008 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_250
timestamp 1663859327
transform 1 0 29344 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_314
timestamp 1663859327
transform 1 0 36512 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_318
timestamp 1663859327
transform 1 0 36960 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_321
timestamp 1663859327
transform 1 0 37296 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_385
timestamp 1663859327
transform 1 0 44464 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_389
timestamp 1663859327
transform 1 0 44912 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_392
timestamp 1663859327
transform 1 0 45248 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_456
timestamp 1663859327
transform 1 0 52416 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_460
timestamp 1663859327
transform 1 0 52864 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_463
timestamp 1663859327
transform 1 0 53200 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_527
timestamp 1663859327
transform 1 0 60368 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_531
timestamp 1663859327
transform 1 0 60816 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_534
timestamp 1663859327
transform 1 0 61152 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_598
timestamp 1663859327
transform 1 0 68320 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_602
timestamp 1663859327
transform 1 0 68768 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_605
timestamp 1663859327
transform 1 0 69104 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_669
timestamp 1663859327
transform 1 0 76272 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_673
timestamp 1663859327
transform 1 0 76720 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_676
timestamp 1663859327
transform 1 0 77056 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_740
timestamp 1663859327
transform 1 0 84224 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_744
timestamp 1663859327
transform 1 0 84672 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_747
timestamp 1663859327
transform 1 0 85008 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_811
timestamp 1663859327
transform 1 0 92176 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_815
timestamp 1663859327
transform 1 0 92624 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_818
timestamp 1663859327
transform 1 0 92960 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_882
timestamp 1663859327
transform 1 0 100128 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_886
timestamp 1663859327
transform 1 0 100576 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_889
timestamp 1663859327
transform 1 0 100912 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_953
timestamp 1663859327
transform 1 0 108080 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_957
timestamp 1663859327
transform 1 0 108528 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_150_960
timestamp 1663859327
transform 1 0 108864 0 1 120736
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_1024
timestamp 1663859327
transform 1 0 116032 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_150_1028
timestamp 1663859327
transform 1 0 116480 0 1 120736
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_150_1031
timestamp 1663859327
transform 1 0 116816 0 1 120736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_150_1039
timestamp 1663859327
transform 1 0 117712 0 1 120736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_150_1043
timestamp 1663859327
transform 1 0 118160 0 1 120736
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_2
timestamp 1663859327
transform 1 0 1568 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_7
timestamp 1663859327
transform 1 0 2128 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_73
timestamp 1663859327
transform 1 0 9520 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_137
timestamp 1663859327
transform 1 0 16688 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_141
timestamp 1663859327
transform 1 0 17136 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_144
timestamp 1663859327
transform 1 0 17472 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_208
timestamp 1663859327
transform 1 0 24640 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_212
timestamp 1663859327
transform 1 0 25088 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_215
timestamp 1663859327
transform 1 0 25424 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_279
timestamp 1663859327
transform 1 0 32592 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_283
timestamp 1663859327
transform 1 0 33040 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_286
timestamp 1663859327
transform 1 0 33376 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_350
timestamp 1663859327
transform 1 0 40544 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_354
timestamp 1663859327
transform 1 0 40992 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_357
timestamp 1663859327
transform 1 0 41328 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_421
timestamp 1663859327
transform 1 0 48496 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_425
timestamp 1663859327
transform 1 0 48944 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_428
timestamp 1663859327
transform 1 0 49280 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_492
timestamp 1663859327
transform 1 0 56448 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_496
timestamp 1663859327
transform 1 0 56896 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_499
timestamp 1663859327
transform 1 0 57232 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_563
timestamp 1663859327
transform 1 0 64400 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_567
timestamp 1663859327
transform 1 0 64848 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_570
timestamp 1663859327
transform 1 0 65184 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_634
timestamp 1663859327
transform 1 0 72352 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_638
timestamp 1663859327
transform 1 0 72800 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_641
timestamp 1663859327
transform 1 0 73136 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_705
timestamp 1663859327
transform 1 0 80304 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_709
timestamp 1663859327
transform 1 0 80752 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_712
timestamp 1663859327
transform 1 0 81088 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_776
timestamp 1663859327
transform 1 0 88256 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_780
timestamp 1663859327
transform 1 0 88704 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_783
timestamp 1663859327
transform 1 0 89040 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_847
timestamp 1663859327
transform 1 0 96208 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_851
timestamp 1663859327
transform 1 0 96656 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_854
timestamp 1663859327
transform 1 0 96992 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_918
timestamp 1663859327
transform 1 0 104160 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_922
timestamp 1663859327
transform 1 0 104608 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_151_925
timestamp 1663859327
transform 1 0 104944 0 -1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_151_989
timestamp 1663859327
transform 1 0 112112 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_993
timestamp 1663859327
transform 1 0 112560 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_151_996
timestamp 1663859327
transform 1 0 112896 0 -1 122304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_151_1028
timestamp 1663859327
transform 1 0 116480 0 -1 122304
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_151_1044
timestamp 1663859327
transform 1 0 118272 0 -1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_152_2
timestamp 1663859327
transform 1 0 1568 0 1 122304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_34
timestamp 1663859327
transform 1 0 5152 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_37
timestamp 1663859327
transform 1 0 5488 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_101
timestamp 1663859327
transform 1 0 12656 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_105
timestamp 1663859327
transform 1 0 13104 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_108
timestamp 1663859327
transform 1 0 13440 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_172
timestamp 1663859327
transform 1 0 20608 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_176
timestamp 1663859327
transform 1 0 21056 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_179
timestamp 1663859327
transform 1 0 21392 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_243
timestamp 1663859327
transform 1 0 28560 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_247
timestamp 1663859327
transform 1 0 29008 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_250
timestamp 1663859327
transform 1 0 29344 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_314
timestamp 1663859327
transform 1 0 36512 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_318
timestamp 1663859327
transform 1 0 36960 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_321
timestamp 1663859327
transform 1 0 37296 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_385
timestamp 1663859327
transform 1 0 44464 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_389
timestamp 1663859327
transform 1 0 44912 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_392
timestamp 1663859327
transform 1 0 45248 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_456
timestamp 1663859327
transform 1 0 52416 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_460
timestamp 1663859327
transform 1 0 52864 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_463
timestamp 1663859327
transform 1 0 53200 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_527
timestamp 1663859327
transform 1 0 60368 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_531
timestamp 1663859327
transform 1 0 60816 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_534
timestamp 1663859327
transform 1 0 61152 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_598
timestamp 1663859327
transform 1 0 68320 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_602
timestamp 1663859327
transform 1 0 68768 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_605
timestamp 1663859327
transform 1 0 69104 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_669
timestamp 1663859327
transform 1 0 76272 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_673
timestamp 1663859327
transform 1 0 76720 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_676
timestamp 1663859327
transform 1 0 77056 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_740
timestamp 1663859327
transform 1 0 84224 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_744
timestamp 1663859327
transform 1 0 84672 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_747
timestamp 1663859327
transform 1 0 85008 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_811
timestamp 1663859327
transform 1 0 92176 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_815
timestamp 1663859327
transform 1 0 92624 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_818
timestamp 1663859327
transform 1 0 92960 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_882
timestamp 1663859327
transform 1 0 100128 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_886
timestamp 1663859327
transform 1 0 100576 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_889
timestamp 1663859327
transform 1 0 100912 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_953
timestamp 1663859327
transform 1 0 108080 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_957
timestamp 1663859327
transform 1 0 108528 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_152_960
timestamp 1663859327
transform 1 0 108864 0 1 122304
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_1024
timestamp 1663859327
transform 1 0 116032 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_152_1028
timestamp 1663859327
transform 1 0 116480 0 1 122304
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_152_1031
timestamp 1663859327
transform 1 0 116816 0 1 122304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_152_1039
timestamp 1663859327
transform 1 0 117712 0 1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_152_1043
timestamp 1663859327
transform 1 0 118160 0 1 122304
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_2
timestamp 1663859327
transform 1 0 1568 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_7
timestamp 1663859327
transform 1 0 2128 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_73
timestamp 1663859327
transform 1 0 9520 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_137
timestamp 1663859327
transform 1 0 16688 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_141
timestamp 1663859327
transform 1 0 17136 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_144
timestamp 1663859327
transform 1 0 17472 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_208
timestamp 1663859327
transform 1 0 24640 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_212
timestamp 1663859327
transform 1 0 25088 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_215
timestamp 1663859327
transform 1 0 25424 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_279
timestamp 1663859327
transform 1 0 32592 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_283
timestamp 1663859327
transform 1 0 33040 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_286
timestamp 1663859327
transform 1 0 33376 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_350
timestamp 1663859327
transform 1 0 40544 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_354
timestamp 1663859327
transform 1 0 40992 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_357
timestamp 1663859327
transform 1 0 41328 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_421
timestamp 1663859327
transform 1 0 48496 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_425
timestamp 1663859327
transform 1 0 48944 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_428
timestamp 1663859327
transform 1 0 49280 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_492
timestamp 1663859327
transform 1 0 56448 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_496
timestamp 1663859327
transform 1 0 56896 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_499
timestamp 1663859327
transform 1 0 57232 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_563
timestamp 1663859327
transform 1 0 64400 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_567
timestamp 1663859327
transform 1 0 64848 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_570
timestamp 1663859327
transform 1 0 65184 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_634
timestamp 1663859327
transform 1 0 72352 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_638
timestamp 1663859327
transform 1 0 72800 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_641
timestamp 1663859327
transform 1 0 73136 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_705
timestamp 1663859327
transform 1 0 80304 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_709
timestamp 1663859327
transform 1 0 80752 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_712
timestamp 1663859327
transform 1 0 81088 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_776
timestamp 1663859327
transform 1 0 88256 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_780
timestamp 1663859327
transform 1 0 88704 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_783
timestamp 1663859327
transform 1 0 89040 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_847
timestamp 1663859327
transform 1 0 96208 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_851
timestamp 1663859327
transform 1 0 96656 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_854
timestamp 1663859327
transform 1 0 96992 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_918
timestamp 1663859327
transform 1 0 104160 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_922
timestamp 1663859327
transform 1 0 104608 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_153_925
timestamp 1663859327
transform 1 0 104944 0 -1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_153_989
timestamp 1663859327
transform 1 0 112112 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_993
timestamp 1663859327
transform 1 0 112560 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_153_996
timestamp 1663859327
transform 1 0 112896 0 -1 123872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_153_1028
timestamp 1663859327
transform 1 0 116480 0 -1 123872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_153_1044
timestamp 1663859327
transform 1 0 118272 0 -1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_154_2
timestamp 1663859327
transform 1 0 1568 0 1 123872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_34
timestamp 1663859327
transform 1 0 5152 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_37
timestamp 1663859327
transform 1 0 5488 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_101
timestamp 1663859327
transform 1 0 12656 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_105
timestamp 1663859327
transform 1 0 13104 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_108
timestamp 1663859327
transform 1 0 13440 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_172
timestamp 1663859327
transform 1 0 20608 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_176
timestamp 1663859327
transform 1 0 21056 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_179
timestamp 1663859327
transform 1 0 21392 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_243
timestamp 1663859327
transform 1 0 28560 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_247
timestamp 1663859327
transform 1 0 29008 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_250
timestamp 1663859327
transform 1 0 29344 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_314
timestamp 1663859327
transform 1 0 36512 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_318
timestamp 1663859327
transform 1 0 36960 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_321
timestamp 1663859327
transform 1 0 37296 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_385
timestamp 1663859327
transform 1 0 44464 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_389
timestamp 1663859327
transform 1 0 44912 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_392
timestamp 1663859327
transform 1 0 45248 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_456
timestamp 1663859327
transform 1 0 52416 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_460
timestamp 1663859327
transform 1 0 52864 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_463
timestamp 1663859327
transform 1 0 53200 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_527
timestamp 1663859327
transform 1 0 60368 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_531
timestamp 1663859327
transform 1 0 60816 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_534
timestamp 1663859327
transform 1 0 61152 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_598
timestamp 1663859327
transform 1 0 68320 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_602
timestamp 1663859327
transform 1 0 68768 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_605
timestamp 1663859327
transform 1 0 69104 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_669
timestamp 1663859327
transform 1 0 76272 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_673
timestamp 1663859327
transform 1 0 76720 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_676
timestamp 1663859327
transform 1 0 77056 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_740
timestamp 1663859327
transform 1 0 84224 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_744
timestamp 1663859327
transform 1 0 84672 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_747
timestamp 1663859327
transform 1 0 85008 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_811
timestamp 1663859327
transform 1 0 92176 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_815
timestamp 1663859327
transform 1 0 92624 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_818
timestamp 1663859327
transform 1 0 92960 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_882
timestamp 1663859327
transform 1 0 100128 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_886
timestamp 1663859327
transform 1 0 100576 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_889
timestamp 1663859327
transform 1 0 100912 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_953
timestamp 1663859327
transform 1 0 108080 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_957
timestamp 1663859327
transform 1 0 108528 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_154_960
timestamp 1663859327
transform 1 0 108864 0 1 123872
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_154_1024
timestamp 1663859327
transform 1 0 116032 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_1028
timestamp 1663859327
transform 1 0 116480 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_154_1031
timestamp 1663859327
transform 1 0 116816 0 1 123872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_1039
timestamp 1663859327
transform 1 0 117712 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_154_1044
timestamp 1663859327
transform 1 0 118272 0 1 123872
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_2
timestamp 1663859327
transform 1 0 1568 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_7
timestamp 1663859327
transform 1 0 2128 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_73
timestamp 1663859327
transform 1 0 9520 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_137
timestamp 1663859327
transform 1 0 16688 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_141
timestamp 1663859327
transform 1 0 17136 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_144
timestamp 1663859327
transform 1 0 17472 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_208
timestamp 1663859327
transform 1 0 24640 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_212
timestamp 1663859327
transform 1 0 25088 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_215
timestamp 1663859327
transform 1 0 25424 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_279
timestamp 1663859327
transform 1 0 32592 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_283
timestamp 1663859327
transform 1 0 33040 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_286
timestamp 1663859327
transform 1 0 33376 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_350
timestamp 1663859327
transform 1 0 40544 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_354
timestamp 1663859327
transform 1 0 40992 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_357
timestamp 1663859327
transform 1 0 41328 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_421
timestamp 1663859327
transform 1 0 48496 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_425
timestamp 1663859327
transform 1 0 48944 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_428
timestamp 1663859327
transform 1 0 49280 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_492
timestamp 1663859327
transform 1 0 56448 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_496
timestamp 1663859327
transform 1 0 56896 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_499
timestamp 1663859327
transform 1 0 57232 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_563
timestamp 1663859327
transform 1 0 64400 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_567
timestamp 1663859327
transform 1 0 64848 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_570
timestamp 1663859327
transform 1 0 65184 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_634
timestamp 1663859327
transform 1 0 72352 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_638
timestamp 1663859327
transform 1 0 72800 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_641
timestamp 1663859327
transform 1 0 73136 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_705
timestamp 1663859327
transform 1 0 80304 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_709
timestamp 1663859327
transform 1 0 80752 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_712
timestamp 1663859327
transform 1 0 81088 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_776
timestamp 1663859327
transform 1 0 88256 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_780
timestamp 1663859327
transform 1 0 88704 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_783
timestamp 1663859327
transform 1 0 89040 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_847
timestamp 1663859327
transform 1 0 96208 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_851
timestamp 1663859327
transform 1 0 96656 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_854
timestamp 1663859327
transform 1 0 96992 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_918
timestamp 1663859327
transform 1 0 104160 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_922
timestamp 1663859327
transform 1 0 104608 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_155_925
timestamp 1663859327
transform 1 0 104944 0 -1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_155_989
timestamp 1663859327
transform 1 0 112112 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_993
timestamp 1663859327
transform 1 0 112560 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_155_996
timestamp 1663859327
transform 1 0 112896 0 -1 125440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_155_1028
timestamp 1663859327
transform 1 0 116480 0 -1 125440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_155_1044
timestamp 1663859327
transform 1 0 118272 0 -1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_156_2
timestamp 1663859327
transform 1 0 1568 0 1 125440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_34
timestamp 1663859327
transform 1 0 5152 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_37
timestamp 1663859327
transform 1 0 5488 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_101
timestamp 1663859327
transform 1 0 12656 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_105
timestamp 1663859327
transform 1 0 13104 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_108
timestamp 1663859327
transform 1 0 13440 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_172
timestamp 1663859327
transform 1 0 20608 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_176
timestamp 1663859327
transform 1 0 21056 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_179
timestamp 1663859327
transform 1 0 21392 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_243
timestamp 1663859327
transform 1 0 28560 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_247
timestamp 1663859327
transform 1 0 29008 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_250
timestamp 1663859327
transform 1 0 29344 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_314
timestamp 1663859327
transform 1 0 36512 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_318
timestamp 1663859327
transform 1 0 36960 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_321
timestamp 1663859327
transform 1 0 37296 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_385
timestamp 1663859327
transform 1 0 44464 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_389
timestamp 1663859327
transform 1 0 44912 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_392
timestamp 1663859327
transform 1 0 45248 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_456
timestamp 1663859327
transform 1 0 52416 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_460
timestamp 1663859327
transform 1 0 52864 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_463
timestamp 1663859327
transform 1 0 53200 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_527
timestamp 1663859327
transform 1 0 60368 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_531
timestamp 1663859327
transform 1 0 60816 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_534
timestamp 1663859327
transform 1 0 61152 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_598
timestamp 1663859327
transform 1 0 68320 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_602
timestamp 1663859327
transform 1 0 68768 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_605
timestamp 1663859327
transform 1 0 69104 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_669
timestamp 1663859327
transform 1 0 76272 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_673
timestamp 1663859327
transform 1 0 76720 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_676
timestamp 1663859327
transform 1 0 77056 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_740
timestamp 1663859327
transform 1 0 84224 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_744
timestamp 1663859327
transform 1 0 84672 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_747
timestamp 1663859327
transform 1 0 85008 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_811
timestamp 1663859327
transform 1 0 92176 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_815
timestamp 1663859327
transform 1 0 92624 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_818
timestamp 1663859327
transform 1 0 92960 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_882
timestamp 1663859327
transform 1 0 100128 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_886
timestamp 1663859327
transform 1 0 100576 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_889
timestamp 1663859327
transform 1 0 100912 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_953
timestamp 1663859327
transform 1 0 108080 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_957
timestamp 1663859327
transform 1 0 108528 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_156_960
timestamp 1663859327
transform 1 0 108864 0 1 125440
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_1024
timestamp 1663859327
transform 1 0 116032 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_156_1028
timestamp 1663859327
transform 1 0 116480 0 1 125440
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_156_1031
timestamp 1663859327
transform 1 0 116816 0 1 125440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_156_1039
timestamp 1663859327
transform 1 0 117712 0 1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_156_1043
timestamp 1663859327
transform 1 0 118160 0 1 125440
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_2
timestamp 1663859327
transform 1 0 1568 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_66
timestamp 1663859327
transform 1 0 8736 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_70
timestamp 1663859327
transform 1 0 9184 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_73
timestamp 1663859327
transform 1 0 9520 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_137
timestamp 1663859327
transform 1 0 16688 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_141
timestamp 1663859327
transform 1 0 17136 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_144
timestamp 1663859327
transform 1 0 17472 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_208
timestamp 1663859327
transform 1 0 24640 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_212
timestamp 1663859327
transform 1 0 25088 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_215
timestamp 1663859327
transform 1 0 25424 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_279
timestamp 1663859327
transform 1 0 32592 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_283
timestamp 1663859327
transform 1 0 33040 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_286
timestamp 1663859327
transform 1 0 33376 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_350
timestamp 1663859327
transform 1 0 40544 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_354
timestamp 1663859327
transform 1 0 40992 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_357
timestamp 1663859327
transform 1 0 41328 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_421
timestamp 1663859327
transform 1 0 48496 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_425
timestamp 1663859327
transform 1 0 48944 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_428
timestamp 1663859327
transform 1 0 49280 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_492
timestamp 1663859327
transform 1 0 56448 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_496
timestamp 1663859327
transform 1 0 56896 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_499
timestamp 1663859327
transform 1 0 57232 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_563
timestamp 1663859327
transform 1 0 64400 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_567
timestamp 1663859327
transform 1 0 64848 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_570
timestamp 1663859327
transform 1 0 65184 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_634
timestamp 1663859327
transform 1 0 72352 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_638
timestamp 1663859327
transform 1 0 72800 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_641
timestamp 1663859327
transform 1 0 73136 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_705
timestamp 1663859327
transform 1 0 80304 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_709
timestamp 1663859327
transform 1 0 80752 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_712
timestamp 1663859327
transform 1 0 81088 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_776
timestamp 1663859327
transform 1 0 88256 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_780
timestamp 1663859327
transform 1 0 88704 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_783
timestamp 1663859327
transform 1 0 89040 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_847
timestamp 1663859327
transform 1 0 96208 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_851
timestamp 1663859327
transform 1 0 96656 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_854
timestamp 1663859327
transform 1 0 96992 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_918
timestamp 1663859327
transform 1 0 104160 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_922
timestamp 1663859327
transform 1 0 104608 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_157_925
timestamp 1663859327
transform 1 0 104944 0 -1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_989
timestamp 1663859327
transform 1 0 112112 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_993
timestamp 1663859327
transform 1 0 112560 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_157_996
timestamp 1663859327
transform 1 0 112896 0 -1 127008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_157_1028
timestamp 1663859327
transform 1 0 116480 0 -1 127008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_157_1036
timestamp 1663859327
transform 1 0 117376 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_157_1044
timestamp 1663859327
transform 1 0 118272 0 -1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_2
timestamp 1663859327
transform 1 0 1568 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_158_7
timestamp 1663859327
transform 1 0 2128 0 1 127008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_158_23
timestamp 1663859327
transform 1 0 3920 0 1 127008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_31
timestamp 1663859327
transform 1 0 4816 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_37
timestamp 1663859327
transform 1 0 5488 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_101
timestamp 1663859327
transform 1 0 12656 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_105
timestamp 1663859327
transform 1 0 13104 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_108
timestamp 1663859327
transform 1 0 13440 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_172
timestamp 1663859327
transform 1 0 20608 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_176
timestamp 1663859327
transform 1 0 21056 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_179
timestamp 1663859327
transform 1 0 21392 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_243
timestamp 1663859327
transform 1 0 28560 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_247
timestamp 1663859327
transform 1 0 29008 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_250
timestamp 1663859327
transform 1 0 29344 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_314
timestamp 1663859327
transform 1 0 36512 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_318
timestamp 1663859327
transform 1 0 36960 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_321
timestamp 1663859327
transform 1 0 37296 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_385
timestamp 1663859327
transform 1 0 44464 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_389
timestamp 1663859327
transform 1 0 44912 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_392
timestamp 1663859327
transform 1 0 45248 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_456
timestamp 1663859327
transform 1 0 52416 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_460
timestamp 1663859327
transform 1 0 52864 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_463
timestamp 1663859327
transform 1 0 53200 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_527
timestamp 1663859327
transform 1 0 60368 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_531
timestamp 1663859327
transform 1 0 60816 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_534
timestamp 1663859327
transform 1 0 61152 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_598
timestamp 1663859327
transform 1 0 68320 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_602
timestamp 1663859327
transform 1 0 68768 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_605
timestamp 1663859327
transform 1 0 69104 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_669
timestamp 1663859327
transform 1 0 76272 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_673
timestamp 1663859327
transform 1 0 76720 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_676
timestamp 1663859327
transform 1 0 77056 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_740
timestamp 1663859327
transform 1 0 84224 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_744
timestamp 1663859327
transform 1 0 84672 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_747
timestamp 1663859327
transform 1 0 85008 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_811
timestamp 1663859327
transform 1 0 92176 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_815
timestamp 1663859327
transform 1 0 92624 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_818
timestamp 1663859327
transform 1 0 92960 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_882
timestamp 1663859327
transform 1 0 100128 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_886
timestamp 1663859327
transform 1 0 100576 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_889
timestamp 1663859327
transform 1 0 100912 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_953
timestamp 1663859327
transform 1 0 108080 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_957
timestamp 1663859327
transform 1 0 108528 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_158_960
timestamp 1663859327
transform 1 0 108864 0 1 127008
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_1024
timestamp 1663859327
transform 1 0 116032 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_158_1028
timestamp 1663859327
transform 1 0 116480 0 1 127008
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_158_1031
timestamp 1663859327
transform 1 0 116816 0 1 127008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_158_1039
timestamp 1663859327
transform 1 0 117712 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_158_1043
timestamp 1663859327
transform 1 0 118160 0 1 127008
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_2
timestamp 1663859327
transform 1 0 1568 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_7
timestamp 1663859327
transform 1 0 2128 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_73
timestamp 1663859327
transform 1 0 9520 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_137
timestamp 1663859327
transform 1 0 16688 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_141
timestamp 1663859327
transform 1 0 17136 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_144
timestamp 1663859327
transform 1 0 17472 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_208
timestamp 1663859327
transform 1 0 24640 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_212
timestamp 1663859327
transform 1 0 25088 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_215
timestamp 1663859327
transform 1 0 25424 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_279
timestamp 1663859327
transform 1 0 32592 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_283
timestamp 1663859327
transform 1 0 33040 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_286
timestamp 1663859327
transform 1 0 33376 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_350
timestamp 1663859327
transform 1 0 40544 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_354
timestamp 1663859327
transform 1 0 40992 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_357
timestamp 1663859327
transform 1 0 41328 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_421
timestamp 1663859327
transform 1 0 48496 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_425
timestamp 1663859327
transform 1 0 48944 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_428
timestamp 1663859327
transform 1 0 49280 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_492
timestamp 1663859327
transform 1 0 56448 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_496
timestamp 1663859327
transform 1 0 56896 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_499
timestamp 1663859327
transform 1 0 57232 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_563
timestamp 1663859327
transform 1 0 64400 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_567
timestamp 1663859327
transform 1 0 64848 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_570
timestamp 1663859327
transform 1 0 65184 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_634
timestamp 1663859327
transform 1 0 72352 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_638
timestamp 1663859327
transform 1 0 72800 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_641
timestamp 1663859327
transform 1 0 73136 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_705
timestamp 1663859327
transform 1 0 80304 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_709
timestamp 1663859327
transform 1 0 80752 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_712
timestamp 1663859327
transform 1 0 81088 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_776
timestamp 1663859327
transform 1 0 88256 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_780
timestamp 1663859327
transform 1 0 88704 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_783
timestamp 1663859327
transform 1 0 89040 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_847
timestamp 1663859327
transform 1 0 96208 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_851
timestamp 1663859327
transform 1 0 96656 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_854
timestamp 1663859327
transform 1 0 96992 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_918
timestamp 1663859327
transform 1 0 104160 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_922
timestamp 1663859327
transform 1 0 104608 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_159_925
timestamp 1663859327
transform 1 0 104944 0 -1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_159_989
timestamp 1663859327
transform 1 0 112112 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_993
timestamp 1663859327
transform 1 0 112560 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_159_996
timestamp 1663859327
transform 1 0 112896 0 -1 128576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_159_1028
timestamp 1663859327
transform 1 0 116480 0 -1 128576
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_159_1044
timestamp 1663859327
transform 1 0 118272 0 -1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_160_2
timestamp 1663859327
transform 1 0 1568 0 1 128576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_34
timestamp 1663859327
transform 1 0 5152 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_37
timestamp 1663859327
transform 1 0 5488 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_101
timestamp 1663859327
transform 1 0 12656 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_105
timestamp 1663859327
transform 1 0 13104 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_108
timestamp 1663859327
transform 1 0 13440 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_172
timestamp 1663859327
transform 1 0 20608 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_176
timestamp 1663859327
transform 1 0 21056 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_179
timestamp 1663859327
transform 1 0 21392 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_243
timestamp 1663859327
transform 1 0 28560 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_247
timestamp 1663859327
transform 1 0 29008 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_250
timestamp 1663859327
transform 1 0 29344 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_314
timestamp 1663859327
transform 1 0 36512 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_318
timestamp 1663859327
transform 1 0 36960 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_321
timestamp 1663859327
transform 1 0 37296 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_385
timestamp 1663859327
transform 1 0 44464 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_389
timestamp 1663859327
transform 1 0 44912 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_392
timestamp 1663859327
transform 1 0 45248 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_456
timestamp 1663859327
transform 1 0 52416 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_460
timestamp 1663859327
transform 1 0 52864 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_463
timestamp 1663859327
transform 1 0 53200 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_527
timestamp 1663859327
transform 1 0 60368 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_531
timestamp 1663859327
transform 1 0 60816 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_534
timestamp 1663859327
transform 1 0 61152 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_598
timestamp 1663859327
transform 1 0 68320 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_602
timestamp 1663859327
transform 1 0 68768 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_605
timestamp 1663859327
transform 1 0 69104 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_669
timestamp 1663859327
transform 1 0 76272 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_673
timestamp 1663859327
transform 1 0 76720 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_676
timestamp 1663859327
transform 1 0 77056 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_740
timestamp 1663859327
transform 1 0 84224 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_744
timestamp 1663859327
transform 1 0 84672 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_747
timestamp 1663859327
transform 1 0 85008 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_811
timestamp 1663859327
transform 1 0 92176 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_815
timestamp 1663859327
transform 1 0 92624 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_818
timestamp 1663859327
transform 1 0 92960 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_882
timestamp 1663859327
transform 1 0 100128 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_886
timestamp 1663859327
transform 1 0 100576 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_889
timestamp 1663859327
transform 1 0 100912 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_953
timestamp 1663859327
transform 1 0 108080 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_957
timestamp 1663859327
transform 1 0 108528 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_160_960
timestamp 1663859327
transform 1 0 108864 0 1 128576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_1024
timestamp 1663859327
transform 1 0 116032 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_160_1028
timestamp 1663859327
transform 1 0 116480 0 1 128576
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_160_1031
timestamp 1663859327
transform 1 0 116816 0 1 128576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_160_1039
timestamp 1663859327
transform 1 0 117712 0 1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_160_1043
timestamp 1663859327
transform 1 0 118160 0 1 128576
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_2
timestamp 1663859327
transform 1 0 1568 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_66
timestamp 1663859327
transform 1 0 8736 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_70
timestamp 1663859327
transform 1 0 9184 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_73
timestamp 1663859327
transform 1 0 9520 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_137
timestamp 1663859327
transform 1 0 16688 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_141
timestamp 1663859327
transform 1 0 17136 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_144
timestamp 1663859327
transform 1 0 17472 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_208
timestamp 1663859327
transform 1 0 24640 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_212
timestamp 1663859327
transform 1 0 25088 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_215
timestamp 1663859327
transform 1 0 25424 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_279
timestamp 1663859327
transform 1 0 32592 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_283
timestamp 1663859327
transform 1 0 33040 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_286
timestamp 1663859327
transform 1 0 33376 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_350
timestamp 1663859327
transform 1 0 40544 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_354
timestamp 1663859327
transform 1 0 40992 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_357
timestamp 1663859327
transform 1 0 41328 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_421
timestamp 1663859327
transform 1 0 48496 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_425
timestamp 1663859327
transform 1 0 48944 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_428
timestamp 1663859327
transform 1 0 49280 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_492
timestamp 1663859327
transform 1 0 56448 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_496
timestamp 1663859327
transform 1 0 56896 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_499
timestamp 1663859327
transform 1 0 57232 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_563
timestamp 1663859327
transform 1 0 64400 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_567
timestamp 1663859327
transform 1 0 64848 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_570
timestamp 1663859327
transform 1 0 65184 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_634
timestamp 1663859327
transform 1 0 72352 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_638
timestamp 1663859327
transform 1 0 72800 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_641
timestamp 1663859327
transform 1 0 73136 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_705
timestamp 1663859327
transform 1 0 80304 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_709
timestamp 1663859327
transform 1 0 80752 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_712
timestamp 1663859327
transform 1 0 81088 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_776
timestamp 1663859327
transform 1 0 88256 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_780
timestamp 1663859327
transform 1 0 88704 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_783
timestamp 1663859327
transform 1 0 89040 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_847
timestamp 1663859327
transform 1 0 96208 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_851
timestamp 1663859327
transform 1 0 96656 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_854
timestamp 1663859327
transform 1 0 96992 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_918
timestamp 1663859327
transform 1 0 104160 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_922
timestamp 1663859327
transform 1 0 104608 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_161_925
timestamp 1663859327
transform 1 0 104944 0 -1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_161_989
timestamp 1663859327
transform 1 0 112112 0 -1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_993
timestamp 1663859327
transform 1 0 112560 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_161_996
timestamp 1663859327
transform 1 0 112896 0 -1 130144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_161_1028
timestamp 1663859327
transform 1 0 116480 0 -1 130144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_161_1044
timestamp 1663859327
transform 1 0 118272 0 -1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_2
timestamp 1663859327
transform 1 0 1568 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_162_7
timestamp 1663859327
transform 1 0 2128 0 1 130144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_162_23
timestamp 1663859327
transform 1 0 3920 0 1 130144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_31
timestamp 1663859327
transform 1 0 4816 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_37
timestamp 1663859327
transform 1 0 5488 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_101
timestamp 1663859327
transform 1 0 12656 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_105
timestamp 1663859327
transform 1 0 13104 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_108
timestamp 1663859327
transform 1 0 13440 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_172
timestamp 1663859327
transform 1 0 20608 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_176
timestamp 1663859327
transform 1 0 21056 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_179
timestamp 1663859327
transform 1 0 21392 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_243
timestamp 1663859327
transform 1 0 28560 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_247
timestamp 1663859327
transform 1 0 29008 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_250
timestamp 1663859327
transform 1 0 29344 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_314
timestamp 1663859327
transform 1 0 36512 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_318
timestamp 1663859327
transform 1 0 36960 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_321
timestamp 1663859327
transform 1 0 37296 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_385
timestamp 1663859327
transform 1 0 44464 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_389
timestamp 1663859327
transform 1 0 44912 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_392
timestamp 1663859327
transform 1 0 45248 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_456
timestamp 1663859327
transform 1 0 52416 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_460
timestamp 1663859327
transform 1 0 52864 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_463
timestamp 1663859327
transform 1 0 53200 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_527
timestamp 1663859327
transform 1 0 60368 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_531
timestamp 1663859327
transform 1 0 60816 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_534
timestamp 1663859327
transform 1 0 61152 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_598
timestamp 1663859327
transform 1 0 68320 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_602
timestamp 1663859327
transform 1 0 68768 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_605
timestamp 1663859327
transform 1 0 69104 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_669
timestamp 1663859327
transform 1 0 76272 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_673
timestamp 1663859327
transform 1 0 76720 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_676
timestamp 1663859327
transform 1 0 77056 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_740
timestamp 1663859327
transform 1 0 84224 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_744
timestamp 1663859327
transform 1 0 84672 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_747
timestamp 1663859327
transform 1 0 85008 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_811
timestamp 1663859327
transform 1 0 92176 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_815
timestamp 1663859327
transform 1 0 92624 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_818
timestamp 1663859327
transform 1 0 92960 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_882
timestamp 1663859327
transform 1 0 100128 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_886
timestamp 1663859327
transform 1 0 100576 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_889
timestamp 1663859327
transform 1 0 100912 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_953
timestamp 1663859327
transform 1 0 108080 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_957
timestamp 1663859327
transform 1 0 108528 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_162_960
timestamp 1663859327
transform 1 0 108864 0 1 130144
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_1024
timestamp 1663859327
transform 1 0 116032 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_162_1028
timestamp 1663859327
transform 1 0 116480 0 1 130144
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_162_1031
timestamp 1663859327
transform 1 0 116816 0 1 130144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_162_1039
timestamp 1663859327
transform 1 0 117712 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_162_1043
timestamp 1663859327
transform 1 0 118160 0 1 130144
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_2
timestamp 1663859327
transform 1 0 1568 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_66
timestamp 1663859327
transform 1 0 8736 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_70
timestamp 1663859327
transform 1 0 9184 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_73
timestamp 1663859327
transform 1 0 9520 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_137
timestamp 1663859327
transform 1 0 16688 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_141
timestamp 1663859327
transform 1 0 17136 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_144
timestamp 1663859327
transform 1 0 17472 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_208
timestamp 1663859327
transform 1 0 24640 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_212
timestamp 1663859327
transform 1 0 25088 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_215
timestamp 1663859327
transform 1 0 25424 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_279
timestamp 1663859327
transform 1 0 32592 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_283
timestamp 1663859327
transform 1 0 33040 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_286
timestamp 1663859327
transform 1 0 33376 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_350
timestamp 1663859327
transform 1 0 40544 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_354
timestamp 1663859327
transform 1 0 40992 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_357
timestamp 1663859327
transform 1 0 41328 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_421
timestamp 1663859327
transform 1 0 48496 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_425
timestamp 1663859327
transform 1 0 48944 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_428
timestamp 1663859327
transform 1 0 49280 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_492
timestamp 1663859327
transform 1 0 56448 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_496
timestamp 1663859327
transform 1 0 56896 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_499
timestamp 1663859327
transform 1 0 57232 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_563
timestamp 1663859327
transform 1 0 64400 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_567
timestamp 1663859327
transform 1 0 64848 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_570
timestamp 1663859327
transform 1 0 65184 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_634
timestamp 1663859327
transform 1 0 72352 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_638
timestamp 1663859327
transform 1 0 72800 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_641
timestamp 1663859327
transform 1 0 73136 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_705
timestamp 1663859327
transform 1 0 80304 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_709
timestamp 1663859327
transform 1 0 80752 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_712
timestamp 1663859327
transform 1 0 81088 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_776
timestamp 1663859327
transform 1 0 88256 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_780
timestamp 1663859327
transform 1 0 88704 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_783
timestamp 1663859327
transform 1 0 89040 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_847
timestamp 1663859327
transform 1 0 96208 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_851
timestamp 1663859327
transform 1 0 96656 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_854
timestamp 1663859327
transform 1 0 96992 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_918
timestamp 1663859327
transform 1 0 104160 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_922
timestamp 1663859327
transform 1 0 104608 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_163_925
timestamp 1663859327
transform 1 0 104944 0 -1 131712
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_163_989
timestamp 1663859327
transform 1 0 112112 0 -1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_993
timestamp 1663859327
transform 1 0 112560 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_163_996
timestamp 1663859327
transform 1 0 112896 0 -1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_163_1028
timestamp 1663859327
transform 1 0 116480 0 -1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_163_1044
timestamp 1663859327
transform 1 0 118272 0 -1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_2
timestamp 1663859327
transform 1 0 1568 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_7
timestamp 1663859327
transform 1 0 2128 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_13
timestamp 1663859327
transform 1 0 2800 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_29
timestamp 1663859327
transform 1 0 4592 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_33
timestamp 1663859327
transform 1 0 5040 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_164_37
timestamp 1663859327
transform 1 0 5488 0 1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_69
timestamp 1663859327
transform 1 0 9072 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_72
timestamp 1663859327
transform 1 0 9408 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_76
timestamp 1663859327
transform 1 0 9856 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_78
timestamp 1663859327
transform 1 0 10080 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_83
timestamp 1663859327
transform 1 0 10640 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_95
timestamp 1663859327
transform 1 0 11984 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_103
timestamp 1663859327
transform 1 0 12880 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_107
timestamp 1663859327
transform 1 0 13328 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_112
timestamp 1663859327
transform 1 0 13888 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_128
timestamp 1663859327
transform 1 0 15680 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_136
timestamp 1663859327
transform 1 0 16576 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_142
timestamp 1663859327
transform 1 0 17248 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_158
timestamp 1663859327
transform 1 0 19040 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_166
timestamp 1663859327
transform 1 0 19936 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_170
timestamp 1663859327
transform 1 0 20384 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_174
timestamp 1663859327
transform 1 0 20832 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_177
timestamp 1663859327
transform 1 0 21168 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_192
timestamp 1663859327
transform 1 0 22848 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_196
timestamp 1663859327
transform 1 0 23296 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_198
timestamp 1663859327
transform 1 0 23520 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_203
timestamp 1663859327
transform 1 0 24080 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_207
timestamp 1663859327
transform 1 0 24528 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_209
timestamp 1663859327
transform 1 0 24752 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_212
timestamp 1663859327
transform 1 0 25088 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_220
timestamp 1663859327
transform 1 0 25984 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_222
timestamp 1663859327
transform 1 0 26208 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_227
timestamp 1663859327
transform 1 0 26768 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_239
timestamp 1663859327
transform 1 0 28112 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_243
timestamp 1663859327
transform 1 0 28560 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_247
timestamp 1663859327
transform 1 0 29008 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_251
timestamp 1663859327
transform 1 0 29456 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_257
timestamp 1663859327
transform 1 0 30128 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_269
timestamp 1663859327
transform 1 0 31472 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_277
timestamp 1663859327
transform 1 0 32368 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_279
timestamp 1663859327
transform 1 0 32592 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_282
timestamp 1663859327
transform 1 0 32928 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_298
timestamp 1663859327
transform 1 0 34720 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_306
timestamp 1663859327
transform 1 0 35616 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_314
timestamp 1663859327
transform 1 0 36512 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_317
timestamp 1663859327
transform 1 0 36848 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_323
timestamp 1663859327
transform 1 0 37520 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_339
timestamp 1663859327
transform 1 0 39312 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_347
timestamp 1663859327
transform 1 0 40208 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_349
timestamp 1663859327
transform 1 0 40432 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_164_352
timestamp 1663859327
transform 1 0 40768 0 1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_384
timestamp 1663859327
transform 1 0 44352 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_387
timestamp 1663859327
transform 1 0 44688 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_395
timestamp 1663859327
transform 1 0 45584 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_401
timestamp 1663859327
transform 1 0 46256 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_417
timestamp 1663859327
transform 1 0 48048 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_419
timestamp 1663859327
transform 1 0 48272 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_422
timestamp 1663859327
transform 1 0 48608 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_438
timestamp 1663859327
transform 1 0 50400 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_442
timestamp 1663859327
transform 1 0 50848 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_444
timestamp 1663859327
transform 1 0 51072 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_449
timestamp 1663859327
transform 1 0 51632 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_453
timestamp 1663859327
transform 1 0 52080 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_457
timestamp 1663859327
transform 1 0 52528 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_461
timestamp 1663859327
transform 1 0 52976 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_467
timestamp 1663859327
transform 1 0 53648 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_479
timestamp 1663859327
transform 1 0 54992 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_487
timestamp 1663859327
transform 1 0 55888 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_489
timestamp 1663859327
transform 1 0 56112 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_492
timestamp 1663859327
transform 1 0 56448 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_508
timestamp 1663859327
transform 1 0 58240 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_510
timestamp 1663859327
transform 1 0 58464 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_515
timestamp 1663859327
transform 1 0 59024 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_519
timestamp 1663859327
transform 1 0 59472 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_521
timestamp 1663859327
transform 1 0 59696 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_524
timestamp 1663859327
transform 1 0 60032 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_527
timestamp 1663859327
transform 1 0 60368 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_534
timestamp 1663859327
transform 1 0 61152 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_540
timestamp 1663859327
transform 1 0 61824 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_548
timestamp 1663859327
transform 1 0 62720 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_552
timestamp 1663859327
transform 1 0 63168 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_557
timestamp 1663859327
transform 1 0 63728 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_559
timestamp 1663859327
transform 1 0 63952 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_562
timestamp 1663859327
transform 1 0 64288 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_564
timestamp 1663859327
transform 1 0 64512 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_569
timestamp 1663859327
transform 1 0 65072 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_581
timestamp 1663859327
transform 1 0 66416 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_593
timestamp 1663859327
transform 1 0 67760 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_597
timestamp 1663859327
transform 1 0 68208 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_605
timestamp 1663859327
transform 1 0 69104 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_611
timestamp 1663859327
transform 1 0 69776 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_627
timestamp 1663859327
transform 1 0 71568 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_629
timestamp 1663859327
transform 1 0 71792 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_632
timestamp 1663859327
transform 1 0 72128 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_637
timestamp 1663859327
transform 1 0 72688 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_641
timestamp 1663859327
transform 1 0 73136 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_647
timestamp 1663859327
transform 1 0 73808 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_659
timestamp 1663859327
transform 1 0 75152 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_663
timestamp 1663859327
transform 1 0 75600 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_667
timestamp 1663859327
transform 1 0 76048 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_672
timestamp 1663859327
transform 1 0 76608 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_688
timestamp 1663859327
transform 1 0 78400 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_696
timestamp 1663859327
transform 1 0 79296 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_702
timestamp 1663859327
transform 1 0 79968 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_706
timestamp 1663859327
transform 1 0 80416 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_708
timestamp 1663859327
transform 1 0 80640 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_713
timestamp 1663859327
transform 1 0 81200 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_725
timestamp 1663859327
transform 1 0 82544 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_733
timestamp 1663859327
transform 1 0 83440 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_737
timestamp 1663859327
transform 1 0 83888 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_743
timestamp 1663859327
transform 1 0 84560 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_755
timestamp 1663859327
transform 1 0 85904 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_763
timestamp 1663859327
transform 1 0 86800 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_767
timestamp 1663859327
transform 1 0 87248 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_769
timestamp 1663859327
transform 1 0 87472 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_772
timestamp 1663859327
transform 1 0 87808 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_774
timestamp 1663859327
transform 1 0 88032 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_779
timestamp 1663859327
transform 1 0 88592 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_791
timestamp 1663859327
transform 1 0 89936 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_799
timestamp 1663859327
transform 1 0 90832 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_803
timestamp 1663859327
transform 1 0 91280 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_164_807
timestamp 1663859327
transform 1 0 91728 0 1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_839
timestamp 1663859327
transform 1 0 95312 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_842
timestamp 1663859327
transform 1 0 95648 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_847
timestamp 1663859327
transform 1 0 96208 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_863
timestamp 1663859327
transform 1 0 98000 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_871
timestamp 1663859327
transform 1 0 98896 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_164_877
timestamp 1663859327
transform 1 0 99568 0 1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_909
timestamp 1663859327
transform 1 0 103152 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_912
timestamp 1663859327
transform 1 0 103488 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_917
timestamp 1663859327
transform 1 0 104048 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_164_923
timestamp 1663859327
transform 1 0 104720 0 1 131712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_939
timestamp 1663859327
transform 1 0 106512 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_943
timestamp 1663859327
transform 1 0 106960 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_947
timestamp 1663859327
transform 1 0 107408 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_955
timestamp 1663859327
transform 1 0 108304 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_959
timestamp 1663859327
transform 1 0 108752 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_164_965
timestamp 1663859327
transform 1 0 109424 0 1 131712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_973
timestamp 1663859327
transform 1 0 110320 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_977
timestamp 1663859327
transform 1 0 110768 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_979
timestamp 1663859327
transform 1 0 110992 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_164_982
timestamp 1663859327
transform 1 0 111328 0 1 131712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_1014
timestamp 1663859327
transform 1 0 114912 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_1017
timestamp 1663859327
transform 1 0 115248 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_164_1022
timestamp 1663859327
transform 1 0 115808 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_164_1026
timestamp 1663859327
transform 1 0 116256 0 1 131712
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_1031
timestamp 1663859327
transform 1 0 116816 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_1037
timestamp 1663859327
transform 1 0 117488 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_164_1043
timestamp 1663859327
transform 1 0 118160 0 1 131712
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1663859327
transform -1 0 118608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1663859327
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1663859327
transform -1 0 118608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1663859327
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1663859327
transform -1 0 118608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1663859327
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1663859327
transform -1 0 118608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1663859327
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1663859327
transform -1 0 118608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1663859327
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1663859327
transform -1 0 118608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1663859327
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1663859327
transform -1 0 118608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1663859327
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1663859327
transform -1 0 118608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1663859327
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1663859327
transform -1 0 118608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1663859327
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1663859327
transform -1 0 118608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1663859327
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1663859327
transform -1 0 118608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1663859327
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1663859327
transform -1 0 118608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1663859327
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1663859327
transform -1 0 118608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1663859327
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1663859327
transform -1 0 118608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1663859327
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1663859327
transform -1 0 118608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1663859327
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1663859327
transform -1 0 118608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1663859327
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1663859327
transform -1 0 118608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1663859327
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1663859327
transform -1 0 118608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1663859327
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1663859327
transform -1 0 118608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1663859327
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1663859327
transform -1 0 118608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1663859327
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1663859327
transform -1 0 118608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1663859327
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1663859327
transform -1 0 118608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1663859327
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1663859327
transform -1 0 118608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1663859327
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1663859327
transform -1 0 118608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1663859327
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1663859327
transform -1 0 118608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1663859327
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1663859327
transform -1 0 118608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1663859327
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1663859327
transform -1 0 118608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1663859327
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1663859327
transform -1 0 118608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1663859327
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1663859327
transform -1 0 118608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1663859327
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1663859327
transform -1 0 118608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1663859327
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1663859327
transform -1 0 118608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1663859327
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1663859327
transform -1 0 118608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1663859327
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1663859327
transform -1 0 118608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1663859327
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1663859327
transform -1 0 118608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1663859327
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1663859327
transform -1 0 118608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1663859327
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1663859327
transform -1 0 118608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1663859327
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1663859327
transform -1 0 118608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1663859327
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1663859327
transform -1 0 118608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1663859327
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1663859327
transform -1 0 118608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1663859327
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1663859327
transform -1 0 118608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1663859327
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1663859327
transform -1 0 118608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1663859327
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1663859327
transform -1 0 118608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1663859327
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1663859327
transform -1 0 118608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1663859327
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1663859327
transform -1 0 118608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1663859327
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1663859327
transform -1 0 118608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1663859327
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1663859327
transform -1 0 118608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1663859327
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1663859327
transform -1 0 118608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1663859327
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1663859327
transform -1 0 118608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1663859327
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1663859327
transform -1 0 118608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1663859327
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1663859327
transform -1 0 118608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1663859327
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1663859327
transform -1 0 118608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1663859327
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1663859327
transform -1 0 118608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1663859327
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1663859327
transform -1 0 118608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1663859327
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1663859327
transform -1 0 118608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1663859327
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1663859327
transform -1 0 118608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1663859327
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1663859327
transform -1 0 118608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1663859327
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1663859327
transform -1 0 118608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1663859327
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1663859327
transform -1 0 118608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1663859327
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1663859327
transform -1 0 118608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1663859327
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1663859327
transform -1 0 118608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1663859327
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1663859327
transform -1 0 118608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1663859327
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1663859327
transform -1 0 118608 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1663859327
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1663859327
transform -1 0 118608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1663859327
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1663859327
transform -1 0 118608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1663859327
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1663859327
transform -1 0 118608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1663859327
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1663859327
transform -1 0 118608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1663859327
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1663859327
transform -1 0 118608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1663859327
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1663859327
transform -1 0 118608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1663859327
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1663859327
transform -1 0 118608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1663859327
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1663859327
transform -1 0 118608 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1663859327
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1663859327
transform -1 0 118608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1663859327
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1663859327
transform -1 0 118608 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1663859327
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1663859327
transform -1 0 118608 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1663859327
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1663859327
transform -1 0 118608 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1663859327
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1663859327
transform -1 0 118608 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1663859327
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1663859327
transform -1 0 118608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1663859327
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1663859327
transform -1 0 118608 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1663859327
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1663859327
transform -1 0 118608 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1663859327
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1663859327
transform -1 0 118608 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1663859327
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1663859327
transform -1 0 118608 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1663859327
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1663859327
transform -1 0 118608 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1663859327
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1663859327
transform -1 0 118608 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1663859327
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1663859327
transform -1 0 118608 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1663859327
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1663859327
transform -1 0 118608 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1663859327
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1663859327
transform -1 0 118608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1663859327
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1663859327
transform -1 0 118608 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1663859327
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1663859327
transform -1 0 118608 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1663859327
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1663859327
transform -1 0 118608 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1663859327
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1663859327
transform -1 0 118608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1663859327
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1663859327
transform -1 0 118608 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1663859327
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1663859327
transform -1 0 118608 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1663859327
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1663859327
transform -1 0 118608 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1663859327
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1663859327
transform -1 0 118608 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1663859327
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1663859327
transform -1 0 118608 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_188
timestamp 1663859327
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_189
timestamp 1663859327
transform -1 0 118608 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_190
timestamp 1663859327
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_191
timestamp 1663859327
transform -1 0 118608 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_192
timestamp 1663859327
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_193
timestamp 1663859327
transform -1 0 118608 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_194
timestamp 1663859327
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_195
timestamp 1663859327
transform -1 0 118608 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_196
timestamp 1663859327
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_197
timestamp 1663859327
transform -1 0 118608 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_198
timestamp 1663859327
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_199
timestamp 1663859327
transform -1 0 118608 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_200
timestamp 1663859327
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_201
timestamp 1663859327
transform -1 0 118608 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_202
timestamp 1663859327
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_203
timestamp 1663859327
transform -1 0 118608 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_204
timestamp 1663859327
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_205
timestamp 1663859327
transform -1 0 118608 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_206
timestamp 1663859327
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_207
timestamp 1663859327
transform -1 0 118608 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_208
timestamp 1663859327
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_209
timestamp 1663859327
transform -1 0 118608 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_210
timestamp 1663859327
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_211
timestamp 1663859327
transform -1 0 118608 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_212
timestamp 1663859327
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_213
timestamp 1663859327
transform -1 0 118608 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_214
timestamp 1663859327
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_215
timestamp 1663859327
transform -1 0 118608 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_216
timestamp 1663859327
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_217
timestamp 1663859327
transform -1 0 118608 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_218
timestamp 1663859327
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_219
timestamp 1663859327
transform -1 0 118608 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_220
timestamp 1663859327
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_221
timestamp 1663859327
transform -1 0 118608 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_222
timestamp 1663859327
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_223
timestamp 1663859327
transform -1 0 118608 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_224
timestamp 1663859327
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_225
timestamp 1663859327
transform -1 0 118608 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_226
timestamp 1663859327
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_227
timestamp 1663859327
transform -1 0 118608 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_228
timestamp 1663859327
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_229
timestamp 1663859327
transform -1 0 118608 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_230
timestamp 1663859327
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_231
timestamp 1663859327
transform -1 0 118608 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_232
timestamp 1663859327
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_233
timestamp 1663859327
transform -1 0 118608 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_234
timestamp 1663859327
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_235
timestamp 1663859327
transform -1 0 118608 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_236
timestamp 1663859327
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_237
timestamp 1663859327
transform -1 0 118608 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_238
timestamp 1663859327
transform 1 0 1344 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_239
timestamp 1663859327
transform -1 0 118608 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_240
timestamp 1663859327
transform 1 0 1344 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_241
timestamp 1663859327
transform -1 0 118608 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_242
timestamp 1663859327
transform 1 0 1344 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_243
timestamp 1663859327
transform -1 0 118608 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_244
timestamp 1663859327
transform 1 0 1344 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_245
timestamp 1663859327
transform -1 0 118608 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_246
timestamp 1663859327
transform 1 0 1344 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_247
timestamp 1663859327
transform -1 0 118608 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_248
timestamp 1663859327
transform 1 0 1344 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_249
timestamp 1663859327
transform -1 0 118608 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_250
timestamp 1663859327
transform 1 0 1344 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_251
timestamp 1663859327
transform -1 0 118608 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_252
timestamp 1663859327
transform 1 0 1344 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_253
timestamp 1663859327
transform -1 0 118608 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_254
timestamp 1663859327
transform 1 0 1344 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_255
timestamp 1663859327
transform -1 0 118608 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_256
timestamp 1663859327
transform 1 0 1344 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_257
timestamp 1663859327
transform -1 0 118608 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_258
timestamp 1663859327
transform 1 0 1344 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_259
timestamp 1663859327
transform -1 0 118608 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_260
timestamp 1663859327
transform 1 0 1344 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_261
timestamp 1663859327
transform -1 0 118608 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_262
timestamp 1663859327
transform 1 0 1344 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_263
timestamp 1663859327
transform -1 0 118608 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_264
timestamp 1663859327
transform 1 0 1344 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_265
timestamp 1663859327
transform -1 0 118608 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_266
timestamp 1663859327
transform 1 0 1344 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_267
timestamp 1663859327
transform -1 0 118608 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_268
timestamp 1663859327
transform 1 0 1344 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_269
timestamp 1663859327
transform -1 0 118608 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_270
timestamp 1663859327
transform 1 0 1344 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_271
timestamp 1663859327
transform -1 0 118608 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_272
timestamp 1663859327
transform 1 0 1344 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_273
timestamp 1663859327
transform -1 0 118608 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_274
timestamp 1663859327
transform 1 0 1344 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_275
timestamp 1663859327
transform -1 0 118608 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_276
timestamp 1663859327
transform 1 0 1344 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_277
timestamp 1663859327
transform -1 0 118608 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_278
timestamp 1663859327
transform 1 0 1344 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_279
timestamp 1663859327
transform -1 0 118608 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_280
timestamp 1663859327
transform 1 0 1344 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_281
timestamp 1663859327
transform -1 0 118608 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_282
timestamp 1663859327
transform 1 0 1344 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_283
timestamp 1663859327
transform -1 0 118608 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_284
timestamp 1663859327
transform 1 0 1344 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_285
timestamp 1663859327
transform -1 0 118608 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_286
timestamp 1663859327
transform 1 0 1344 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_287
timestamp 1663859327
transform -1 0 118608 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_288
timestamp 1663859327
transform 1 0 1344 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_289
timestamp 1663859327
transform -1 0 118608 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_290
timestamp 1663859327
transform 1 0 1344 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_291
timestamp 1663859327
transform -1 0 118608 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_292
timestamp 1663859327
transform 1 0 1344 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_293
timestamp 1663859327
transform -1 0 118608 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_294
timestamp 1663859327
transform 1 0 1344 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_295
timestamp 1663859327
transform -1 0 118608 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_296
timestamp 1663859327
transform 1 0 1344 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_297
timestamp 1663859327
transform -1 0 118608 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_298
timestamp 1663859327
transform 1 0 1344 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_299
timestamp 1663859327
transform -1 0 118608 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_300
timestamp 1663859327
transform 1 0 1344 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_301
timestamp 1663859327
transform -1 0 118608 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_302
timestamp 1663859327
transform 1 0 1344 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_303
timestamp 1663859327
transform -1 0 118608 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_304
timestamp 1663859327
transform 1 0 1344 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_305
timestamp 1663859327
transform -1 0 118608 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_306
timestamp 1663859327
transform 1 0 1344 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_307
timestamp 1663859327
transform -1 0 118608 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_308
timestamp 1663859327
transform 1 0 1344 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_309
timestamp 1663859327
transform -1 0 118608 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_310
timestamp 1663859327
transform 1 0 1344 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_311
timestamp 1663859327
transform -1 0 118608 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_312
timestamp 1663859327
transform 1 0 1344 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_313
timestamp 1663859327
transform -1 0 118608 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_314
timestamp 1663859327
transform 1 0 1344 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_315
timestamp 1663859327
transform -1 0 118608 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_316
timestamp 1663859327
transform 1 0 1344 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_317
timestamp 1663859327
transform -1 0 118608 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_318
timestamp 1663859327
transform 1 0 1344 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_319
timestamp 1663859327
transform -1 0 118608 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_320
timestamp 1663859327
transform 1 0 1344 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_321
timestamp 1663859327
transform -1 0 118608 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_322
timestamp 1663859327
transform 1 0 1344 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_323
timestamp 1663859327
transform -1 0 118608 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_324
timestamp 1663859327
transform 1 0 1344 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_325
timestamp 1663859327
transform -1 0 118608 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_326
timestamp 1663859327
transform 1 0 1344 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_327
timestamp 1663859327
transform -1 0 118608 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_328
timestamp 1663859327
transform 1 0 1344 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_329
timestamp 1663859327
transform -1 0 118608 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1663859327
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1663859327
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1663859327
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1663859327
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1663859327
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1663859327
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1663859327
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1663859327
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1663859327
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1663859327
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1663859327
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1663859327
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1663859327
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1663859327
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1663859327
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1663859327
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1663859327
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1663859327
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1663859327
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1663859327
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1663859327
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1663859327
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1663859327
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1663859327
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1663859327
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1663859327
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1663859327
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1663859327
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1663859327
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1663859327
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1663859327
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1663859327
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1663859327
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1663859327
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1663859327
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1663859327
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1663859327
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1663859327
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1663859327
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1663859327
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1663859327
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1663859327
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1663859327
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1663859327
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1663859327
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1663859327
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1663859327
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1663859327
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1663859327
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1663859327
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1663859327
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1663859327
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1663859327
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1663859327
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1663859327
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1663859327
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1663859327
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1663859327
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1663859327
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1663859327
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1663859327
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1663859327
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1663859327
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1663859327
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1663859327
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1663859327
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1663859327
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1663859327
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1663859327
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1663859327
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1663859327
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1663859327
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1663859327
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1663859327
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1663859327
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1663859327
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1663859327
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1663859327
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1663859327
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1663859327
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1663859327
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1663859327
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1663859327
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1663859327
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1663859327
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1663859327
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1663859327
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1663859327
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1663859327
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1663859327
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1663859327
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1663859327
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1663859327
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1663859327
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1663859327
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1663859327
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1663859327
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1663859327
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1663859327
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1663859327
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1663859327
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1663859327
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1663859327
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1663859327
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1663859327
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1663859327
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1663859327
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1663859327
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1663859327
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1663859327
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1663859327
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1663859327
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1663859327
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1663859327
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1663859327
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1663859327
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1663859327
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1663859327
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1663859327
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1663859327
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1663859327
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1663859327
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1663859327
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1663859327
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1663859327
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1663859327
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1663859327
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1663859327
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1663859327
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1663859327
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1663859327
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1663859327
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1663859327
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1663859327
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1663859327
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1663859327
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1663859327
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1663859327
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1663859327
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1663859327
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1663859327
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1663859327
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1663859327
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1663859327
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1663859327
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1663859327
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1663859327
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1663859327
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1663859327
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1663859327
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1663859327
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1663859327
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1663859327
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1663859327
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1663859327
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1663859327
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1663859327
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1663859327
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1663859327
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1663859327
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1663859327
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1663859327
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1663859327
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1663859327
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1663859327
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1663859327
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1663859327
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1663859327
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1663859327
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1663859327
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1663859327
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1663859327
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1663859327
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1663859327
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1663859327
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1663859327
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1663859327
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1663859327
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1663859327
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1663859327
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1663859327
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1663859327
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1663859327
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1663859327
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1663859327
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1663859327
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1663859327
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1663859327
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1663859327
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1663859327
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1663859327
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1663859327
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1663859327
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1663859327
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1663859327
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1663859327
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1663859327
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1663859327
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1663859327
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1663859327
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1663859327
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1663859327
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1663859327
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1663859327
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1663859327
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1663859327
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1663859327
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1663859327
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1663859327
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1663859327
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1663859327
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1663859327
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1663859327
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1663859327
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1663859327
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1663859327
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1663859327
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1663859327
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1663859327
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1663859327
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1663859327
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1663859327
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1663859327
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1663859327
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1663859327
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1663859327
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1663859327
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1663859327
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1663859327
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1663859327
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1663859327
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1663859327
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1663859327
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1663859327
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1663859327
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1663859327
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1663859327
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1663859327
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1663859327
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1663859327
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1663859327
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1663859327
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1663859327
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1663859327
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1663859327
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1663859327
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1663859327
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1663859327
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1663859327
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1663859327
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1663859327
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1663859327
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1663859327
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1663859327
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1663859327
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1663859327
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1663859327
transform 1 0 92736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1663859327
transform 1 0 100688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1663859327
transform 1 0 108640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1663859327
transform 1 0 116592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1663859327
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1663859327
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1663859327
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1663859327
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1663859327
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1663859327
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1663859327
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1663859327
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1663859327
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1663859327
transform 1 0 80864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1663859327
transform 1 0 88816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1663859327
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1663859327
transform 1 0 104720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1663859327
transform 1 0 112672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1663859327
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1663859327
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1663859327
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1663859327
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1663859327
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1663859327
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1663859327
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1663859327
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1663859327
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1663859327
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1663859327
transform 1 0 84784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1663859327
transform 1 0 92736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1663859327
transform 1 0 100688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1663859327
transform 1 0 108640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1663859327
transform 1 0 116592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1663859327
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1663859327
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1663859327
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1663859327
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1663859327
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1663859327
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1663859327
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1663859327
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1663859327
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1663859327
transform 1 0 80864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1663859327
transform 1 0 88816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1663859327
transform 1 0 96768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1663859327
transform 1 0 104720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1663859327
transform 1 0 112672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1663859327
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1663859327
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1663859327
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1663859327
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1663859327
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1663859327
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1663859327
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1663859327
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1663859327
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1663859327
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1663859327
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1663859327
transform 1 0 92736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1663859327
transform 1 0 100688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1663859327
transform 1 0 108640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1663859327
transform 1 0 116592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1663859327
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1663859327
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1663859327
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1663859327
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1663859327
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1663859327
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1663859327
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1663859327
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1663859327
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1663859327
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1663859327
transform 1 0 88816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1663859327
transform 1 0 96768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1663859327
transform 1 0 104720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1663859327
transform 1 0 112672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1663859327
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1663859327
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1663859327
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1663859327
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1663859327
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1663859327
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1663859327
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1663859327
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1663859327
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1663859327
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1663859327
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1663859327
transform 1 0 92736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1663859327
transform 1 0 100688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1663859327
transform 1 0 108640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1663859327
transform 1 0 116592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1663859327
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1663859327
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1663859327
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1663859327
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1663859327
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1663859327
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1663859327
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1663859327
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1663859327
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1663859327
transform 1 0 80864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1663859327
transform 1 0 88816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1663859327
transform 1 0 96768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1663859327
transform 1 0 104720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1663859327
transform 1 0 112672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1663859327
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1663859327
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1663859327
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1663859327
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1663859327
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1663859327
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1663859327
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1663859327
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1663859327
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1663859327
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1663859327
transform 1 0 84784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1663859327
transform 1 0 92736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1663859327
transform 1 0 100688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1663859327
transform 1 0 108640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1663859327
transform 1 0 116592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1663859327
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1663859327
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1663859327
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1663859327
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1663859327
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1663859327
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1663859327
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1663859327
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1663859327
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1663859327
transform 1 0 80864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1663859327
transform 1 0 88816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1663859327
transform 1 0 96768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1663859327
transform 1 0 104720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1663859327
transform 1 0 112672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1663859327
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1663859327
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1663859327
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1663859327
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1663859327
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1663859327
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1663859327
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1663859327
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1663859327
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1663859327
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1663859327
transform 1 0 84784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1663859327
transform 1 0 92736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1663859327
transform 1 0 100688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1663859327
transform 1 0 108640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1663859327
transform 1 0 116592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1663859327
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1663859327
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1663859327
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1663859327
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1663859327
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1663859327
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1663859327
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1663859327
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1663859327
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1663859327
transform 1 0 80864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1663859327
transform 1 0 88816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1663859327
transform 1 0 96768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1663859327
transform 1 0 104720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1663859327
transform 1 0 112672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1663859327
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1663859327
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1663859327
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1663859327
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1663859327
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1663859327
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1663859327
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1663859327
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1663859327
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1663859327
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1663859327
transform 1 0 84784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1663859327
transform 1 0 92736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1663859327
transform 1 0 100688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1663859327
transform 1 0 108640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1663859327
transform 1 0 116592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1663859327
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1663859327
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1663859327
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1663859327
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1663859327
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1663859327
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1663859327
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1663859327
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1663859327
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1663859327
transform 1 0 80864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1663859327
transform 1 0 88816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1663859327
transform 1 0 96768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1663859327
transform 1 0 104720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1663859327
transform 1 0 112672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1663859327
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1663859327
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1663859327
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1663859327
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1663859327
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1663859327
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1663859327
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1663859327
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1663859327
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1663859327
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1663859327
transform 1 0 84784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1663859327
transform 1 0 92736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1663859327
transform 1 0 100688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1663859327
transform 1 0 108640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1663859327
transform 1 0 116592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1663859327
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1663859327
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1663859327
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1663859327
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1663859327
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1663859327
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1663859327
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1663859327
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1663859327
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1663859327
transform 1 0 80864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1663859327
transform 1 0 88816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1663859327
transform 1 0 96768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1663859327
transform 1 0 104720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1663859327
transform 1 0 112672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1663859327
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1663859327
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1663859327
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1663859327
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1663859327
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1663859327
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1663859327
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1663859327
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1663859327
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1663859327
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1663859327
transform 1 0 84784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1663859327
transform 1 0 92736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1663859327
transform 1 0 100688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1663859327
transform 1 0 108640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1663859327
transform 1 0 116592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1663859327
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1663859327
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1663859327
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1663859327
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1663859327
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1663859327
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1663859327
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1663859327
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1663859327
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1663859327
transform 1 0 80864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1663859327
transform 1 0 88816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1663859327
transform 1 0 96768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1663859327
transform 1 0 104720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1663859327
transform 1 0 112672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1663859327
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1663859327
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1663859327
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1663859327
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1663859327
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1663859327
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1663859327
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1663859327
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1663859327
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1663859327
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1663859327
transform 1 0 84784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1663859327
transform 1 0 92736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1663859327
transform 1 0 100688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1663859327
transform 1 0 108640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1663859327
transform 1 0 116592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1663859327
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1663859327
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1663859327
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1663859327
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1663859327
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1663859327
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1663859327
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1663859327
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1663859327
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1663859327
transform 1 0 80864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1663859327
transform 1 0 88816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1663859327
transform 1 0 96768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1663859327
transform 1 0 104720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1663859327
transform 1 0 112672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1663859327
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1663859327
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1663859327
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1663859327
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1663859327
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1663859327
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1663859327
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1663859327
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1663859327
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1663859327
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1663859327
transform 1 0 84784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1663859327
transform 1 0 92736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1663859327
transform 1 0 100688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1663859327
transform 1 0 108640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1663859327
transform 1 0 116592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1663859327
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1663859327
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1663859327
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1663859327
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1663859327
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1663859327
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1663859327
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1663859327
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1663859327
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1663859327
transform 1 0 80864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1663859327
transform 1 0 88816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1663859327
transform 1 0 96768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1663859327
transform 1 0 104720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1663859327
transform 1 0 112672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1663859327
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1663859327
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1663859327
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_898
timestamp 1663859327
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_899
timestamp 1663859327
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_900
timestamp 1663859327
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_901
timestamp 1663859327
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_902
timestamp 1663859327
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_903
timestamp 1663859327
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_904
timestamp 1663859327
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_905
timestamp 1663859327
transform 1 0 84784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_906
timestamp 1663859327
transform 1 0 92736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_907
timestamp 1663859327
transform 1 0 100688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_908
timestamp 1663859327
transform 1 0 108640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_909
timestamp 1663859327
transform 1 0 116592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_910
timestamp 1663859327
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_911
timestamp 1663859327
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_912
timestamp 1663859327
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_913
timestamp 1663859327
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_914
timestamp 1663859327
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_915
timestamp 1663859327
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_916
timestamp 1663859327
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_917
timestamp 1663859327
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_918
timestamp 1663859327
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_919
timestamp 1663859327
transform 1 0 80864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_920
timestamp 1663859327
transform 1 0 88816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_921
timestamp 1663859327
transform 1 0 96768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_922
timestamp 1663859327
transform 1 0 104720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_923
timestamp 1663859327
transform 1 0 112672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_924
timestamp 1663859327
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_925
timestamp 1663859327
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_926
timestamp 1663859327
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_927
timestamp 1663859327
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_928
timestamp 1663859327
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_929
timestamp 1663859327
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_930
timestamp 1663859327
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_931
timestamp 1663859327
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_932
timestamp 1663859327
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_933
timestamp 1663859327
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_934
timestamp 1663859327
transform 1 0 84784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_935
timestamp 1663859327
transform 1 0 92736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_936
timestamp 1663859327
transform 1 0 100688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_937
timestamp 1663859327
transform 1 0 108640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_938
timestamp 1663859327
transform 1 0 116592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_939
timestamp 1663859327
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_940
timestamp 1663859327
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_941
timestamp 1663859327
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_942
timestamp 1663859327
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_943
timestamp 1663859327
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_944
timestamp 1663859327
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_945
timestamp 1663859327
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_946
timestamp 1663859327
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_947
timestamp 1663859327
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_948
timestamp 1663859327
transform 1 0 80864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_949
timestamp 1663859327
transform 1 0 88816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_950
timestamp 1663859327
transform 1 0 96768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_951
timestamp 1663859327
transform 1 0 104720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_952
timestamp 1663859327
transform 1 0 112672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_953
timestamp 1663859327
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_954
timestamp 1663859327
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_955
timestamp 1663859327
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_956
timestamp 1663859327
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_957
timestamp 1663859327
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_958
timestamp 1663859327
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_959
timestamp 1663859327
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_960
timestamp 1663859327
transform 1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_961
timestamp 1663859327
transform 1 0 68880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_962
timestamp 1663859327
transform 1 0 76832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_963
timestamp 1663859327
transform 1 0 84784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_964
timestamp 1663859327
transform 1 0 92736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_965
timestamp 1663859327
transform 1 0 100688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_966
timestamp 1663859327
transform 1 0 108640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_967
timestamp 1663859327
transform 1 0 116592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_968
timestamp 1663859327
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_969
timestamp 1663859327
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_970
timestamp 1663859327
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_971
timestamp 1663859327
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_972
timestamp 1663859327
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_973
timestamp 1663859327
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_974
timestamp 1663859327
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_975
timestamp 1663859327
transform 1 0 64960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_976
timestamp 1663859327
transform 1 0 72912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_977
timestamp 1663859327
transform 1 0 80864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_978
timestamp 1663859327
transform 1 0 88816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_979
timestamp 1663859327
transform 1 0 96768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_980
timestamp 1663859327
transform 1 0 104720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_981
timestamp 1663859327
transform 1 0 112672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_982
timestamp 1663859327
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_983
timestamp 1663859327
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_984
timestamp 1663859327
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_985
timestamp 1663859327
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_986
timestamp 1663859327
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_987
timestamp 1663859327
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_988
timestamp 1663859327
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_989
timestamp 1663859327
transform 1 0 60928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_990
timestamp 1663859327
transform 1 0 68880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_991
timestamp 1663859327
transform 1 0 76832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_992
timestamp 1663859327
transform 1 0 84784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_993
timestamp 1663859327
transform 1 0 92736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_994
timestamp 1663859327
transform 1 0 100688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_995
timestamp 1663859327
transform 1 0 108640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_996
timestamp 1663859327
transform 1 0 116592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_997
timestamp 1663859327
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_998
timestamp 1663859327
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_999
timestamp 1663859327
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1000
timestamp 1663859327
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1001
timestamp 1663859327
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1002
timestamp 1663859327
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1003
timestamp 1663859327
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1004
timestamp 1663859327
transform 1 0 64960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1005
timestamp 1663859327
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1006
timestamp 1663859327
transform 1 0 80864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1007
timestamp 1663859327
transform 1 0 88816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1008
timestamp 1663859327
transform 1 0 96768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1009
timestamp 1663859327
transform 1 0 104720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1010
timestamp 1663859327
transform 1 0 112672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1011
timestamp 1663859327
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1012
timestamp 1663859327
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1013
timestamp 1663859327
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1014
timestamp 1663859327
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1015
timestamp 1663859327
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1016
timestamp 1663859327
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1017
timestamp 1663859327
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1018
timestamp 1663859327
transform 1 0 60928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1019
timestamp 1663859327
transform 1 0 68880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1020
timestamp 1663859327
transform 1 0 76832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1021
timestamp 1663859327
transform 1 0 84784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1022
timestamp 1663859327
transform 1 0 92736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1023
timestamp 1663859327
transform 1 0 100688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1024
timestamp 1663859327
transform 1 0 108640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1025
timestamp 1663859327
transform 1 0 116592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1026
timestamp 1663859327
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1027
timestamp 1663859327
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1028
timestamp 1663859327
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1029
timestamp 1663859327
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1030
timestamp 1663859327
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1031
timestamp 1663859327
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1032
timestamp 1663859327
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1033
timestamp 1663859327
transform 1 0 64960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1034
timestamp 1663859327
transform 1 0 72912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1035
timestamp 1663859327
transform 1 0 80864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1036
timestamp 1663859327
transform 1 0 88816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1037
timestamp 1663859327
transform 1 0 96768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1038
timestamp 1663859327
transform 1 0 104720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1039
timestamp 1663859327
transform 1 0 112672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1040
timestamp 1663859327
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1041
timestamp 1663859327
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1042
timestamp 1663859327
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1043
timestamp 1663859327
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1044
timestamp 1663859327
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1045
timestamp 1663859327
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1046
timestamp 1663859327
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1047
timestamp 1663859327
transform 1 0 60928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1048
timestamp 1663859327
transform 1 0 68880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1049
timestamp 1663859327
transform 1 0 76832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1050
timestamp 1663859327
transform 1 0 84784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1051
timestamp 1663859327
transform 1 0 92736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1052
timestamp 1663859327
transform 1 0 100688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1053
timestamp 1663859327
transform 1 0 108640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1054
timestamp 1663859327
transform 1 0 116592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1055
timestamp 1663859327
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1056
timestamp 1663859327
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1057
timestamp 1663859327
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1058
timestamp 1663859327
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1059
timestamp 1663859327
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1060
timestamp 1663859327
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1061
timestamp 1663859327
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1062
timestamp 1663859327
transform 1 0 64960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1063
timestamp 1663859327
transform 1 0 72912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1064
timestamp 1663859327
transform 1 0 80864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1065
timestamp 1663859327
transform 1 0 88816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1066
timestamp 1663859327
transform 1 0 96768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1067
timestamp 1663859327
transform 1 0 104720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1068
timestamp 1663859327
transform 1 0 112672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1069
timestamp 1663859327
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1070
timestamp 1663859327
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1071
timestamp 1663859327
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1072
timestamp 1663859327
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1073
timestamp 1663859327
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1074
timestamp 1663859327
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1075
timestamp 1663859327
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1076
timestamp 1663859327
transform 1 0 60928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1077
timestamp 1663859327
transform 1 0 68880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1078
timestamp 1663859327
transform 1 0 76832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1079
timestamp 1663859327
transform 1 0 84784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1080
timestamp 1663859327
transform 1 0 92736 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1081
timestamp 1663859327
transform 1 0 100688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1082
timestamp 1663859327
transform 1 0 108640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1083
timestamp 1663859327
transform 1 0 116592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1084
timestamp 1663859327
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1085
timestamp 1663859327
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1086
timestamp 1663859327
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1087
timestamp 1663859327
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1088
timestamp 1663859327
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1089
timestamp 1663859327
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1090
timestamp 1663859327
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1091
timestamp 1663859327
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1092
timestamp 1663859327
transform 1 0 72912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1093
timestamp 1663859327
transform 1 0 80864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1094
timestamp 1663859327
transform 1 0 88816 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1095
timestamp 1663859327
transform 1 0 96768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1096
timestamp 1663859327
transform 1 0 104720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1097
timestamp 1663859327
transform 1 0 112672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1098
timestamp 1663859327
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1099
timestamp 1663859327
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1100
timestamp 1663859327
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1101
timestamp 1663859327
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1102
timestamp 1663859327
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1103
timestamp 1663859327
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1104
timestamp 1663859327
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1105
timestamp 1663859327
transform 1 0 60928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1106
timestamp 1663859327
transform 1 0 68880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1107
timestamp 1663859327
transform 1 0 76832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1108
timestamp 1663859327
transform 1 0 84784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1109
timestamp 1663859327
transform 1 0 92736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1110
timestamp 1663859327
transform 1 0 100688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1111
timestamp 1663859327
transform 1 0 108640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1112
timestamp 1663859327
transform 1 0 116592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1113
timestamp 1663859327
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1114
timestamp 1663859327
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1115
timestamp 1663859327
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1116
timestamp 1663859327
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1117
timestamp 1663859327
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1118
timestamp 1663859327
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1119
timestamp 1663859327
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1120
timestamp 1663859327
transform 1 0 64960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1121
timestamp 1663859327
transform 1 0 72912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1122
timestamp 1663859327
transform 1 0 80864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1123
timestamp 1663859327
transform 1 0 88816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1124
timestamp 1663859327
transform 1 0 96768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1125
timestamp 1663859327
transform 1 0 104720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1126
timestamp 1663859327
transform 1 0 112672 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1127
timestamp 1663859327
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1128
timestamp 1663859327
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1129
timestamp 1663859327
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1130
timestamp 1663859327
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1131
timestamp 1663859327
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1132
timestamp 1663859327
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1133
timestamp 1663859327
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1134
timestamp 1663859327
transform 1 0 60928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1135
timestamp 1663859327
transform 1 0 68880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1136
timestamp 1663859327
transform 1 0 76832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1137
timestamp 1663859327
transform 1 0 84784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1138
timestamp 1663859327
transform 1 0 92736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1139
timestamp 1663859327
transform 1 0 100688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1140
timestamp 1663859327
transform 1 0 108640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1141
timestamp 1663859327
transform 1 0 116592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1142
timestamp 1663859327
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1143
timestamp 1663859327
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1144
timestamp 1663859327
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1145
timestamp 1663859327
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1146
timestamp 1663859327
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1147
timestamp 1663859327
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1148
timestamp 1663859327
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1149
timestamp 1663859327
transform 1 0 64960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1150
timestamp 1663859327
transform 1 0 72912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1151
timestamp 1663859327
transform 1 0 80864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1152
timestamp 1663859327
transform 1 0 88816 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1153
timestamp 1663859327
transform 1 0 96768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1154
timestamp 1663859327
transform 1 0 104720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1155
timestamp 1663859327
transform 1 0 112672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1156
timestamp 1663859327
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1157
timestamp 1663859327
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1158
timestamp 1663859327
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1159
timestamp 1663859327
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1160
timestamp 1663859327
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1161
timestamp 1663859327
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1162
timestamp 1663859327
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1163
timestamp 1663859327
transform 1 0 60928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1164
timestamp 1663859327
transform 1 0 68880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1165
timestamp 1663859327
transform 1 0 76832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1166
timestamp 1663859327
transform 1 0 84784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1167
timestamp 1663859327
transform 1 0 92736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1168
timestamp 1663859327
transform 1 0 100688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1169
timestamp 1663859327
transform 1 0 108640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1170
timestamp 1663859327
transform 1 0 116592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1171
timestamp 1663859327
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1172
timestamp 1663859327
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1173
timestamp 1663859327
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1174
timestamp 1663859327
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1175
timestamp 1663859327
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1176
timestamp 1663859327
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1177
timestamp 1663859327
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1178
timestamp 1663859327
transform 1 0 64960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1179
timestamp 1663859327
transform 1 0 72912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1180
timestamp 1663859327
transform 1 0 80864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1181
timestamp 1663859327
transform 1 0 88816 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1182
timestamp 1663859327
transform 1 0 96768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1183
timestamp 1663859327
transform 1 0 104720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1184
timestamp 1663859327
transform 1 0 112672 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1185
timestamp 1663859327
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1186
timestamp 1663859327
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1187
timestamp 1663859327
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1188
timestamp 1663859327
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1189
timestamp 1663859327
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1190
timestamp 1663859327
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1191
timestamp 1663859327
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1192
timestamp 1663859327
transform 1 0 60928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1193
timestamp 1663859327
transform 1 0 68880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1194
timestamp 1663859327
transform 1 0 76832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1195
timestamp 1663859327
transform 1 0 84784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1196
timestamp 1663859327
transform 1 0 92736 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1197
timestamp 1663859327
transform 1 0 100688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1198
timestamp 1663859327
transform 1 0 108640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1199
timestamp 1663859327
transform 1 0 116592 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1200
timestamp 1663859327
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1201
timestamp 1663859327
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1202
timestamp 1663859327
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1203
timestamp 1663859327
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1204
timestamp 1663859327
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1205
timestamp 1663859327
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1206
timestamp 1663859327
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1207
timestamp 1663859327
transform 1 0 64960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1208
timestamp 1663859327
transform 1 0 72912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1209
timestamp 1663859327
transform 1 0 80864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1210
timestamp 1663859327
transform 1 0 88816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1211
timestamp 1663859327
transform 1 0 96768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1212
timestamp 1663859327
transform 1 0 104720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1213
timestamp 1663859327
transform 1 0 112672 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1214
timestamp 1663859327
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1215
timestamp 1663859327
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1216
timestamp 1663859327
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1217
timestamp 1663859327
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1218
timestamp 1663859327
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1219
timestamp 1663859327
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1220
timestamp 1663859327
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1221
timestamp 1663859327
transform 1 0 60928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1222
timestamp 1663859327
transform 1 0 68880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1223
timestamp 1663859327
transform 1 0 76832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1224
timestamp 1663859327
transform 1 0 84784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1225
timestamp 1663859327
transform 1 0 92736 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1226
timestamp 1663859327
transform 1 0 100688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1227
timestamp 1663859327
transform 1 0 108640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1228
timestamp 1663859327
transform 1 0 116592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1229
timestamp 1663859327
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1230
timestamp 1663859327
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1231
timestamp 1663859327
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1232
timestamp 1663859327
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1233
timestamp 1663859327
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1234
timestamp 1663859327
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1235
timestamp 1663859327
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1236
timestamp 1663859327
transform 1 0 64960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1237
timestamp 1663859327
transform 1 0 72912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1238
timestamp 1663859327
transform 1 0 80864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1239
timestamp 1663859327
transform 1 0 88816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1240
timestamp 1663859327
transform 1 0 96768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1241
timestamp 1663859327
transform 1 0 104720 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1242
timestamp 1663859327
transform 1 0 112672 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1243
timestamp 1663859327
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1244
timestamp 1663859327
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1245
timestamp 1663859327
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1246
timestamp 1663859327
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1247
timestamp 1663859327
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1248
timestamp 1663859327
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1249
timestamp 1663859327
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1250
timestamp 1663859327
transform 1 0 60928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1251
timestamp 1663859327
transform 1 0 68880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1252
timestamp 1663859327
transform 1 0 76832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1253
timestamp 1663859327
transform 1 0 84784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1254
timestamp 1663859327
transform 1 0 92736 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1255
timestamp 1663859327
transform 1 0 100688 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1256
timestamp 1663859327
transform 1 0 108640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1257
timestamp 1663859327
transform 1 0 116592 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1258
timestamp 1663859327
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1259
timestamp 1663859327
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1260
timestamp 1663859327
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1261
timestamp 1663859327
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1262
timestamp 1663859327
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1263
timestamp 1663859327
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1264
timestamp 1663859327
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1265
timestamp 1663859327
transform 1 0 64960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1266
timestamp 1663859327
transform 1 0 72912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1267
timestamp 1663859327
transform 1 0 80864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1268
timestamp 1663859327
transform 1 0 88816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1269
timestamp 1663859327
transform 1 0 96768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1270
timestamp 1663859327
transform 1 0 104720 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1271
timestamp 1663859327
transform 1 0 112672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1272
timestamp 1663859327
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1273
timestamp 1663859327
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1274
timestamp 1663859327
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1275
timestamp 1663859327
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1276
timestamp 1663859327
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1277
timestamp 1663859327
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1278
timestamp 1663859327
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1279
timestamp 1663859327
transform 1 0 60928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1280
timestamp 1663859327
transform 1 0 68880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1281
timestamp 1663859327
transform 1 0 76832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1282
timestamp 1663859327
transform 1 0 84784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1283
timestamp 1663859327
transform 1 0 92736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1284
timestamp 1663859327
transform 1 0 100688 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1285
timestamp 1663859327
transform 1 0 108640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1286
timestamp 1663859327
transform 1 0 116592 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1287
timestamp 1663859327
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1288
timestamp 1663859327
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1289
timestamp 1663859327
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1290
timestamp 1663859327
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1291
timestamp 1663859327
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1292
timestamp 1663859327
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1293
timestamp 1663859327
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1294
timestamp 1663859327
transform 1 0 64960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1295
timestamp 1663859327
transform 1 0 72912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1296
timestamp 1663859327
transform 1 0 80864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1297
timestamp 1663859327
transform 1 0 88816 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1298
timestamp 1663859327
transform 1 0 96768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1299
timestamp 1663859327
transform 1 0 104720 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1300
timestamp 1663859327
transform 1 0 112672 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1301
timestamp 1663859327
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1302
timestamp 1663859327
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1303
timestamp 1663859327
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1304
timestamp 1663859327
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1305
timestamp 1663859327
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1306
timestamp 1663859327
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1307
timestamp 1663859327
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1308
timestamp 1663859327
transform 1 0 60928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1309
timestamp 1663859327
transform 1 0 68880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1310
timestamp 1663859327
transform 1 0 76832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1311
timestamp 1663859327
transform 1 0 84784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1312
timestamp 1663859327
transform 1 0 92736 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1313
timestamp 1663859327
transform 1 0 100688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1314
timestamp 1663859327
transform 1 0 108640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1315
timestamp 1663859327
transform 1 0 116592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1316
timestamp 1663859327
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1317
timestamp 1663859327
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1318
timestamp 1663859327
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1319
timestamp 1663859327
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1320
timestamp 1663859327
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1321
timestamp 1663859327
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1322
timestamp 1663859327
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1323
timestamp 1663859327
transform 1 0 64960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1324
timestamp 1663859327
transform 1 0 72912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1325
timestamp 1663859327
transform 1 0 80864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1326
timestamp 1663859327
transform 1 0 88816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1327
timestamp 1663859327
transform 1 0 96768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1328
timestamp 1663859327
transform 1 0 104720 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1329
timestamp 1663859327
transform 1 0 112672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1330
timestamp 1663859327
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1331
timestamp 1663859327
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1332
timestamp 1663859327
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1333
timestamp 1663859327
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1334
timestamp 1663859327
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1335
timestamp 1663859327
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1336
timestamp 1663859327
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1337
timestamp 1663859327
transform 1 0 60928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1338
timestamp 1663859327
transform 1 0 68880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1339
timestamp 1663859327
transform 1 0 76832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1340
timestamp 1663859327
transform 1 0 84784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1341
timestamp 1663859327
transform 1 0 92736 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1342
timestamp 1663859327
transform 1 0 100688 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1343
timestamp 1663859327
transform 1 0 108640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1344
timestamp 1663859327
transform 1 0 116592 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1345
timestamp 1663859327
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1346
timestamp 1663859327
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1347
timestamp 1663859327
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1348
timestamp 1663859327
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1349
timestamp 1663859327
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1350
timestamp 1663859327
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1351
timestamp 1663859327
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1352
timestamp 1663859327
transform 1 0 64960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1353
timestamp 1663859327
transform 1 0 72912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1354
timestamp 1663859327
transform 1 0 80864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1355
timestamp 1663859327
transform 1 0 88816 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1356
timestamp 1663859327
transform 1 0 96768 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1357
timestamp 1663859327
transform 1 0 104720 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1358
timestamp 1663859327
transform 1 0 112672 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1359
timestamp 1663859327
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1360
timestamp 1663859327
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1361
timestamp 1663859327
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1362
timestamp 1663859327
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1363
timestamp 1663859327
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1364
timestamp 1663859327
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1365
timestamp 1663859327
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1366
timestamp 1663859327
transform 1 0 60928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1367
timestamp 1663859327
transform 1 0 68880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1368
timestamp 1663859327
transform 1 0 76832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1369
timestamp 1663859327
transform 1 0 84784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1370
timestamp 1663859327
transform 1 0 92736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1371
timestamp 1663859327
transform 1 0 100688 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1372
timestamp 1663859327
transform 1 0 108640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1373
timestamp 1663859327
transform 1 0 116592 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1374
timestamp 1663859327
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1375
timestamp 1663859327
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1376
timestamp 1663859327
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1377
timestamp 1663859327
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1378
timestamp 1663859327
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1379
timestamp 1663859327
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1380
timestamp 1663859327
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1381
timestamp 1663859327
transform 1 0 64960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1382
timestamp 1663859327
transform 1 0 72912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1383
timestamp 1663859327
transform 1 0 80864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1384
timestamp 1663859327
transform 1 0 88816 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1385
timestamp 1663859327
transform 1 0 96768 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1386
timestamp 1663859327
transform 1 0 104720 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1387
timestamp 1663859327
transform 1 0 112672 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1388
timestamp 1663859327
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1389
timestamp 1663859327
transform 1 0 13216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1390
timestamp 1663859327
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1391
timestamp 1663859327
transform 1 0 29120 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1392
timestamp 1663859327
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1393
timestamp 1663859327
transform 1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1394
timestamp 1663859327
transform 1 0 52976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1395
timestamp 1663859327
transform 1 0 60928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1396
timestamp 1663859327
transform 1 0 68880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1397
timestamp 1663859327
transform 1 0 76832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1398
timestamp 1663859327
transform 1 0 84784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1399
timestamp 1663859327
transform 1 0 92736 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1400
timestamp 1663859327
transform 1 0 100688 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1401
timestamp 1663859327
transform 1 0 108640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1402
timestamp 1663859327
transform 1 0 116592 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1403
timestamp 1663859327
transform 1 0 9296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1404
timestamp 1663859327
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1405
timestamp 1663859327
transform 1 0 25200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1406
timestamp 1663859327
transform 1 0 33152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1407
timestamp 1663859327
transform 1 0 41104 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1408
timestamp 1663859327
transform 1 0 49056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1409
timestamp 1663859327
transform 1 0 57008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1410
timestamp 1663859327
transform 1 0 64960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1411
timestamp 1663859327
transform 1 0 72912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1412
timestamp 1663859327
transform 1 0 80864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1413
timestamp 1663859327
transform 1 0 88816 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1414
timestamp 1663859327
transform 1 0 96768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1415
timestamp 1663859327
transform 1 0 104720 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1416
timestamp 1663859327
transform 1 0 112672 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1417
timestamp 1663859327
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1418
timestamp 1663859327
transform 1 0 13216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1419
timestamp 1663859327
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1420
timestamp 1663859327
transform 1 0 29120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1421
timestamp 1663859327
transform 1 0 37072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1422
timestamp 1663859327
transform 1 0 45024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1423
timestamp 1663859327
transform 1 0 52976 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1424
timestamp 1663859327
transform 1 0 60928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1425
timestamp 1663859327
transform 1 0 68880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1426
timestamp 1663859327
transform 1 0 76832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1427
timestamp 1663859327
transform 1 0 84784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1428
timestamp 1663859327
transform 1 0 92736 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1429
timestamp 1663859327
transform 1 0 100688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1430
timestamp 1663859327
transform 1 0 108640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1431
timestamp 1663859327
transform 1 0 116592 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1432
timestamp 1663859327
transform 1 0 9296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1433
timestamp 1663859327
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1434
timestamp 1663859327
transform 1 0 25200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1435
timestamp 1663859327
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1436
timestamp 1663859327
transform 1 0 41104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1437
timestamp 1663859327
transform 1 0 49056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1438
timestamp 1663859327
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1439
timestamp 1663859327
transform 1 0 64960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1440
timestamp 1663859327
transform 1 0 72912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1441
timestamp 1663859327
transform 1 0 80864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1442
timestamp 1663859327
transform 1 0 88816 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1443
timestamp 1663859327
transform 1 0 96768 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1444
timestamp 1663859327
transform 1 0 104720 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1445
timestamp 1663859327
transform 1 0 112672 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1446
timestamp 1663859327
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1447
timestamp 1663859327
transform 1 0 13216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1448
timestamp 1663859327
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1449
timestamp 1663859327
transform 1 0 29120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1450
timestamp 1663859327
transform 1 0 37072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1451
timestamp 1663859327
transform 1 0 45024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1452
timestamp 1663859327
transform 1 0 52976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1453
timestamp 1663859327
transform 1 0 60928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1454
timestamp 1663859327
transform 1 0 68880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1455
timestamp 1663859327
transform 1 0 76832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1456
timestamp 1663859327
transform 1 0 84784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1457
timestamp 1663859327
transform 1 0 92736 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1458
timestamp 1663859327
transform 1 0 100688 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1459
timestamp 1663859327
transform 1 0 108640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1460
timestamp 1663859327
transform 1 0 116592 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1461
timestamp 1663859327
transform 1 0 9296 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1462
timestamp 1663859327
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1463
timestamp 1663859327
transform 1 0 25200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1464
timestamp 1663859327
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1465
timestamp 1663859327
transform 1 0 41104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1466
timestamp 1663859327
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1467
timestamp 1663859327
transform 1 0 57008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1468
timestamp 1663859327
transform 1 0 64960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1469
timestamp 1663859327
transform 1 0 72912 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1470
timestamp 1663859327
transform 1 0 80864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1471
timestamp 1663859327
transform 1 0 88816 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1472
timestamp 1663859327
transform 1 0 96768 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1473
timestamp 1663859327
transform 1 0 104720 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1474
timestamp 1663859327
transform 1 0 112672 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1475
timestamp 1663859327
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1476
timestamp 1663859327
transform 1 0 13216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1477
timestamp 1663859327
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1478
timestamp 1663859327
transform 1 0 29120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1479
timestamp 1663859327
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1480
timestamp 1663859327
transform 1 0 45024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1481
timestamp 1663859327
transform 1 0 52976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1482
timestamp 1663859327
transform 1 0 60928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1483
timestamp 1663859327
transform 1 0 68880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1484
timestamp 1663859327
transform 1 0 76832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1485
timestamp 1663859327
transform 1 0 84784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1486
timestamp 1663859327
transform 1 0 92736 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1487
timestamp 1663859327
transform 1 0 100688 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1488
timestamp 1663859327
transform 1 0 108640 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1489
timestamp 1663859327
transform 1 0 116592 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1490
timestamp 1663859327
transform 1 0 9296 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1491
timestamp 1663859327
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1492
timestamp 1663859327
transform 1 0 25200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1493
timestamp 1663859327
transform 1 0 33152 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1494
timestamp 1663859327
transform 1 0 41104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1495
timestamp 1663859327
transform 1 0 49056 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1496
timestamp 1663859327
transform 1 0 57008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1497
timestamp 1663859327
transform 1 0 64960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1498
timestamp 1663859327
transform 1 0 72912 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1499
timestamp 1663859327
transform 1 0 80864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1500
timestamp 1663859327
transform 1 0 88816 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1501
timestamp 1663859327
transform 1 0 96768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1502
timestamp 1663859327
transform 1 0 104720 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1503
timestamp 1663859327
transform 1 0 112672 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1504
timestamp 1663859327
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1505
timestamp 1663859327
transform 1 0 13216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1506
timestamp 1663859327
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1507
timestamp 1663859327
transform 1 0 29120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1508
timestamp 1663859327
transform 1 0 37072 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1509
timestamp 1663859327
transform 1 0 45024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1510
timestamp 1663859327
transform 1 0 52976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1511
timestamp 1663859327
transform 1 0 60928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1512
timestamp 1663859327
transform 1 0 68880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1513
timestamp 1663859327
transform 1 0 76832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1514
timestamp 1663859327
transform 1 0 84784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1515
timestamp 1663859327
transform 1 0 92736 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1516
timestamp 1663859327
transform 1 0 100688 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1517
timestamp 1663859327
transform 1 0 108640 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1518
timestamp 1663859327
transform 1 0 116592 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1519
timestamp 1663859327
transform 1 0 9296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1520
timestamp 1663859327
transform 1 0 17248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1521
timestamp 1663859327
transform 1 0 25200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1522
timestamp 1663859327
transform 1 0 33152 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1523
timestamp 1663859327
transform 1 0 41104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1524
timestamp 1663859327
transform 1 0 49056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1525
timestamp 1663859327
transform 1 0 57008 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1526
timestamp 1663859327
transform 1 0 64960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1527
timestamp 1663859327
transform 1 0 72912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1528
timestamp 1663859327
transform 1 0 80864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1529
timestamp 1663859327
transform 1 0 88816 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1530
timestamp 1663859327
transform 1 0 96768 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1531
timestamp 1663859327
transform 1 0 104720 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1532
timestamp 1663859327
transform 1 0 112672 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1533
timestamp 1663859327
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1534
timestamp 1663859327
transform 1 0 13216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1535
timestamp 1663859327
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1536
timestamp 1663859327
transform 1 0 29120 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1537
timestamp 1663859327
transform 1 0 37072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1538
timestamp 1663859327
transform 1 0 45024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1539
timestamp 1663859327
transform 1 0 52976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1540
timestamp 1663859327
transform 1 0 60928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1541
timestamp 1663859327
transform 1 0 68880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1542
timestamp 1663859327
transform 1 0 76832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1543
timestamp 1663859327
transform 1 0 84784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1544
timestamp 1663859327
transform 1 0 92736 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1545
timestamp 1663859327
transform 1 0 100688 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1546
timestamp 1663859327
transform 1 0 108640 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1547
timestamp 1663859327
transform 1 0 116592 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1548
timestamp 1663859327
transform 1 0 9296 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1549
timestamp 1663859327
transform 1 0 17248 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1550
timestamp 1663859327
transform 1 0 25200 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1551
timestamp 1663859327
transform 1 0 33152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1552
timestamp 1663859327
transform 1 0 41104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1553
timestamp 1663859327
transform 1 0 49056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1554
timestamp 1663859327
transform 1 0 57008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1555
timestamp 1663859327
transform 1 0 64960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1556
timestamp 1663859327
transform 1 0 72912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1557
timestamp 1663859327
transform 1 0 80864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1558
timestamp 1663859327
transform 1 0 88816 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1559
timestamp 1663859327
transform 1 0 96768 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1560
timestamp 1663859327
transform 1 0 104720 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1561
timestamp 1663859327
transform 1 0 112672 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1562
timestamp 1663859327
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1563
timestamp 1663859327
transform 1 0 13216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1564
timestamp 1663859327
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1565
timestamp 1663859327
transform 1 0 29120 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1566
timestamp 1663859327
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1567
timestamp 1663859327
transform 1 0 45024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1568
timestamp 1663859327
transform 1 0 52976 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1569
timestamp 1663859327
transform 1 0 60928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1570
timestamp 1663859327
transform 1 0 68880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1571
timestamp 1663859327
transform 1 0 76832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1572
timestamp 1663859327
transform 1 0 84784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1573
timestamp 1663859327
transform 1 0 92736 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1574
timestamp 1663859327
transform 1 0 100688 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1575
timestamp 1663859327
transform 1 0 108640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1576
timestamp 1663859327
transform 1 0 116592 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1577
timestamp 1663859327
transform 1 0 9296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1578
timestamp 1663859327
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1579
timestamp 1663859327
transform 1 0 25200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1580
timestamp 1663859327
transform 1 0 33152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1581
timestamp 1663859327
transform 1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1582
timestamp 1663859327
transform 1 0 49056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1583
timestamp 1663859327
transform 1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1584
timestamp 1663859327
transform 1 0 64960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1585
timestamp 1663859327
transform 1 0 72912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1586
timestamp 1663859327
transform 1 0 80864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1587
timestamp 1663859327
transform 1 0 88816 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1588
timestamp 1663859327
transform 1 0 96768 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1589
timestamp 1663859327
transform 1 0 104720 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1590
timestamp 1663859327
transform 1 0 112672 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1591
timestamp 1663859327
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1592
timestamp 1663859327
transform 1 0 13216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1593
timestamp 1663859327
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1594
timestamp 1663859327
transform 1 0 29120 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1595
timestamp 1663859327
transform 1 0 37072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1596
timestamp 1663859327
transform 1 0 45024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1597
timestamp 1663859327
transform 1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1598
timestamp 1663859327
transform 1 0 60928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1599
timestamp 1663859327
transform 1 0 68880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1600
timestamp 1663859327
transform 1 0 76832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1601
timestamp 1663859327
transform 1 0 84784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1602
timestamp 1663859327
transform 1 0 92736 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1603
timestamp 1663859327
transform 1 0 100688 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1604
timestamp 1663859327
transform 1 0 108640 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1605
timestamp 1663859327
transform 1 0 116592 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1606
timestamp 1663859327
transform 1 0 9296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1607
timestamp 1663859327
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1608
timestamp 1663859327
transform 1 0 25200 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1609
timestamp 1663859327
transform 1 0 33152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1610
timestamp 1663859327
transform 1 0 41104 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1611
timestamp 1663859327
transform 1 0 49056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1612
timestamp 1663859327
transform 1 0 57008 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1613
timestamp 1663859327
transform 1 0 64960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1614
timestamp 1663859327
transform 1 0 72912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1615
timestamp 1663859327
transform 1 0 80864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1616
timestamp 1663859327
transform 1 0 88816 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1617
timestamp 1663859327
transform 1 0 96768 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1618
timestamp 1663859327
transform 1 0 104720 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1619
timestamp 1663859327
transform 1 0 112672 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1620
timestamp 1663859327
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1621
timestamp 1663859327
transform 1 0 13216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1622
timestamp 1663859327
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1623
timestamp 1663859327
transform 1 0 29120 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1624
timestamp 1663859327
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1625
timestamp 1663859327
transform 1 0 45024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1626
timestamp 1663859327
transform 1 0 52976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1627
timestamp 1663859327
transform 1 0 60928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1628
timestamp 1663859327
transform 1 0 68880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1629
timestamp 1663859327
transform 1 0 76832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1630
timestamp 1663859327
transform 1 0 84784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1631
timestamp 1663859327
transform 1 0 92736 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1632
timestamp 1663859327
transform 1 0 100688 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1633
timestamp 1663859327
transform 1 0 108640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1634
timestamp 1663859327
transform 1 0 116592 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1635
timestamp 1663859327
transform 1 0 9296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1636
timestamp 1663859327
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1637
timestamp 1663859327
transform 1 0 25200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1638
timestamp 1663859327
transform 1 0 33152 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1639
timestamp 1663859327
transform 1 0 41104 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1640
timestamp 1663859327
transform 1 0 49056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1641
timestamp 1663859327
transform 1 0 57008 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1642
timestamp 1663859327
transform 1 0 64960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1643
timestamp 1663859327
transform 1 0 72912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1644
timestamp 1663859327
transform 1 0 80864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1645
timestamp 1663859327
transform 1 0 88816 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1646
timestamp 1663859327
transform 1 0 96768 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1647
timestamp 1663859327
transform 1 0 104720 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1648
timestamp 1663859327
transform 1 0 112672 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1649
timestamp 1663859327
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1650
timestamp 1663859327
transform 1 0 13216 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1651
timestamp 1663859327
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1652
timestamp 1663859327
transform 1 0 29120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1653
timestamp 1663859327
transform 1 0 37072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1654
timestamp 1663859327
transform 1 0 45024 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1655
timestamp 1663859327
transform 1 0 52976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1656
timestamp 1663859327
transform 1 0 60928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1657
timestamp 1663859327
transform 1 0 68880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1658
timestamp 1663859327
transform 1 0 76832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1659
timestamp 1663859327
transform 1 0 84784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1660
timestamp 1663859327
transform 1 0 92736 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1661
timestamp 1663859327
transform 1 0 100688 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1662
timestamp 1663859327
transform 1 0 108640 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1663
timestamp 1663859327
transform 1 0 116592 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1664
timestamp 1663859327
transform 1 0 9296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1665
timestamp 1663859327
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1666
timestamp 1663859327
transform 1 0 25200 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1667
timestamp 1663859327
transform 1 0 33152 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1668
timestamp 1663859327
transform 1 0 41104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1669
timestamp 1663859327
transform 1 0 49056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1670
timestamp 1663859327
transform 1 0 57008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1671
timestamp 1663859327
transform 1 0 64960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1672
timestamp 1663859327
transform 1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1673
timestamp 1663859327
transform 1 0 80864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1674
timestamp 1663859327
transform 1 0 88816 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1675
timestamp 1663859327
transform 1 0 96768 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1676
timestamp 1663859327
transform 1 0 104720 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1677
timestamp 1663859327
transform 1 0 112672 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1678
timestamp 1663859327
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1679
timestamp 1663859327
transform 1 0 13216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1680
timestamp 1663859327
transform 1 0 21168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1681
timestamp 1663859327
transform 1 0 29120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1682
timestamp 1663859327
transform 1 0 37072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1683
timestamp 1663859327
transform 1 0 45024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1684
timestamp 1663859327
transform 1 0 52976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1685
timestamp 1663859327
transform 1 0 60928 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1686
timestamp 1663859327
transform 1 0 68880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1687
timestamp 1663859327
transform 1 0 76832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1688
timestamp 1663859327
transform 1 0 84784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1689
timestamp 1663859327
transform 1 0 92736 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1690
timestamp 1663859327
transform 1 0 100688 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1691
timestamp 1663859327
transform 1 0 108640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1692
timestamp 1663859327
transform 1 0 116592 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1693
timestamp 1663859327
transform 1 0 9296 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1694
timestamp 1663859327
transform 1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1695
timestamp 1663859327
transform 1 0 25200 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1696
timestamp 1663859327
transform 1 0 33152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1697
timestamp 1663859327
transform 1 0 41104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1698
timestamp 1663859327
transform 1 0 49056 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1699
timestamp 1663859327
transform 1 0 57008 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1700
timestamp 1663859327
transform 1 0 64960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1701
timestamp 1663859327
transform 1 0 72912 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1702
timestamp 1663859327
transform 1 0 80864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1703
timestamp 1663859327
transform 1 0 88816 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1704
timestamp 1663859327
transform 1 0 96768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1705
timestamp 1663859327
transform 1 0 104720 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1706
timestamp 1663859327
transform 1 0 112672 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1707
timestamp 1663859327
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1708
timestamp 1663859327
transform 1 0 13216 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1709
timestamp 1663859327
transform 1 0 21168 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1710
timestamp 1663859327
transform 1 0 29120 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1711
timestamp 1663859327
transform 1 0 37072 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1712
timestamp 1663859327
transform 1 0 45024 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1713
timestamp 1663859327
transform 1 0 52976 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1714
timestamp 1663859327
transform 1 0 60928 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1715
timestamp 1663859327
transform 1 0 68880 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1716
timestamp 1663859327
transform 1 0 76832 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1717
timestamp 1663859327
transform 1 0 84784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1718
timestamp 1663859327
transform 1 0 92736 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1719
timestamp 1663859327
transform 1 0 100688 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1720
timestamp 1663859327
transform 1 0 108640 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1721
timestamp 1663859327
transform 1 0 116592 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1722
timestamp 1663859327
transform 1 0 9296 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1723
timestamp 1663859327
transform 1 0 17248 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1724
timestamp 1663859327
transform 1 0 25200 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1725
timestamp 1663859327
transform 1 0 33152 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1726
timestamp 1663859327
transform 1 0 41104 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1727
timestamp 1663859327
transform 1 0 49056 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1728
timestamp 1663859327
transform 1 0 57008 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1729
timestamp 1663859327
transform 1 0 64960 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1730
timestamp 1663859327
transform 1 0 72912 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1731
timestamp 1663859327
transform 1 0 80864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1732
timestamp 1663859327
transform 1 0 88816 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1733
timestamp 1663859327
transform 1 0 96768 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1734
timestamp 1663859327
transform 1 0 104720 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1735
timestamp 1663859327
transform 1 0 112672 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1736
timestamp 1663859327
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1737
timestamp 1663859327
transform 1 0 13216 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1738
timestamp 1663859327
transform 1 0 21168 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1739
timestamp 1663859327
transform 1 0 29120 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1740
timestamp 1663859327
transform 1 0 37072 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1741
timestamp 1663859327
transform 1 0 45024 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1742
timestamp 1663859327
transform 1 0 52976 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1743
timestamp 1663859327
transform 1 0 60928 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1744
timestamp 1663859327
transform 1 0 68880 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1745
timestamp 1663859327
transform 1 0 76832 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1746
timestamp 1663859327
transform 1 0 84784 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1747
timestamp 1663859327
transform 1 0 92736 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1748
timestamp 1663859327
transform 1 0 100688 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1749
timestamp 1663859327
transform 1 0 108640 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1750
timestamp 1663859327
transform 1 0 116592 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1751
timestamp 1663859327
transform 1 0 9296 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1752
timestamp 1663859327
transform 1 0 17248 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1753
timestamp 1663859327
transform 1 0 25200 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1754
timestamp 1663859327
transform 1 0 33152 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1755
timestamp 1663859327
transform 1 0 41104 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1756
timestamp 1663859327
transform 1 0 49056 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1757
timestamp 1663859327
transform 1 0 57008 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1758
timestamp 1663859327
transform 1 0 64960 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1759
timestamp 1663859327
transform 1 0 72912 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1760
timestamp 1663859327
transform 1 0 80864 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1761
timestamp 1663859327
transform 1 0 88816 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1762
timestamp 1663859327
transform 1 0 96768 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1763
timestamp 1663859327
transform 1 0 104720 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1764
timestamp 1663859327
transform 1 0 112672 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1765
timestamp 1663859327
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1766
timestamp 1663859327
transform 1 0 13216 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1767
timestamp 1663859327
transform 1 0 21168 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1768
timestamp 1663859327
transform 1 0 29120 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1769
timestamp 1663859327
transform 1 0 37072 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1770
timestamp 1663859327
transform 1 0 45024 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1771
timestamp 1663859327
transform 1 0 52976 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1772
timestamp 1663859327
transform 1 0 60928 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1773
timestamp 1663859327
transform 1 0 68880 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1774
timestamp 1663859327
transform 1 0 76832 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1775
timestamp 1663859327
transform 1 0 84784 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1776
timestamp 1663859327
transform 1 0 92736 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1777
timestamp 1663859327
transform 1 0 100688 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1778
timestamp 1663859327
transform 1 0 108640 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1779
timestamp 1663859327
transform 1 0 116592 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1780
timestamp 1663859327
transform 1 0 9296 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1781
timestamp 1663859327
transform 1 0 17248 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1782
timestamp 1663859327
transform 1 0 25200 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1783
timestamp 1663859327
transform 1 0 33152 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1784
timestamp 1663859327
transform 1 0 41104 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1785
timestamp 1663859327
transform 1 0 49056 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1786
timestamp 1663859327
transform 1 0 57008 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1787
timestamp 1663859327
transform 1 0 64960 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1788
timestamp 1663859327
transform 1 0 72912 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1789
timestamp 1663859327
transform 1 0 80864 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1790
timestamp 1663859327
transform 1 0 88816 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1791
timestamp 1663859327
transform 1 0 96768 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1792
timestamp 1663859327
transform 1 0 104720 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1793
timestamp 1663859327
transform 1 0 112672 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1794
timestamp 1663859327
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1795
timestamp 1663859327
transform 1 0 13216 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1796
timestamp 1663859327
transform 1 0 21168 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1797
timestamp 1663859327
transform 1 0 29120 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1798
timestamp 1663859327
transform 1 0 37072 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1799
timestamp 1663859327
transform 1 0 45024 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1800
timestamp 1663859327
transform 1 0 52976 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1801
timestamp 1663859327
transform 1 0 60928 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1802
timestamp 1663859327
transform 1 0 68880 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1803
timestamp 1663859327
transform 1 0 76832 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1804
timestamp 1663859327
transform 1 0 84784 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1805
timestamp 1663859327
transform 1 0 92736 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1806
timestamp 1663859327
transform 1 0 100688 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1807
timestamp 1663859327
transform 1 0 108640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1808
timestamp 1663859327
transform 1 0 116592 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1809
timestamp 1663859327
transform 1 0 9296 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1810
timestamp 1663859327
transform 1 0 17248 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1811
timestamp 1663859327
transform 1 0 25200 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1812
timestamp 1663859327
transform 1 0 33152 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1813
timestamp 1663859327
transform 1 0 41104 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1814
timestamp 1663859327
transform 1 0 49056 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1815
timestamp 1663859327
transform 1 0 57008 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1816
timestamp 1663859327
transform 1 0 64960 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1817
timestamp 1663859327
transform 1 0 72912 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1818
timestamp 1663859327
transform 1 0 80864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1819
timestamp 1663859327
transform 1 0 88816 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1820
timestamp 1663859327
transform 1 0 96768 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1821
timestamp 1663859327
transform 1 0 104720 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1822
timestamp 1663859327
transform 1 0 112672 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1823
timestamp 1663859327
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1824
timestamp 1663859327
transform 1 0 13216 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1825
timestamp 1663859327
transform 1 0 21168 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1826
timestamp 1663859327
transform 1 0 29120 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1827
timestamp 1663859327
transform 1 0 37072 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1828
timestamp 1663859327
transform 1 0 45024 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1829
timestamp 1663859327
transform 1 0 52976 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1830
timestamp 1663859327
transform 1 0 60928 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1831
timestamp 1663859327
transform 1 0 68880 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1832
timestamp 1663859327
transform 1 0 76832 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1833
timestamp 1663859327
transform 1 0 84784 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1834
timestamp 1663859327
transform 1 0 92736 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1835
timestamp 1663859327
transform 1 0 100688 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1836
timestamp 1663859327
transform 1 0 108640 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1837
timestamp 1663859327
transform 1 0 116592 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1838
timestamp 1663859327
transform 1 0 9296 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1839
timestamp 1663859327
transform 1 0 17248 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1840
timestamp 1663859327
transform 1 0 25200 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1841
timestamp 1663859327
transform 1 0 33152 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1842
timestamp 1663859327
transform 1 0 41104 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1843
timestamp 1663859327
transform 1 0 49056 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1844
timestamp 1663859327
transform 1 0 57008 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1845
timestamp 1663859327
transform 1 0 64960 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1846
timestamp 1663859327
transform 1 0 72912 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1847
timestamp 1663859327
transform 1 0 80864 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1848
timestamp 1663859327
transform 1 0 88816 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1849
timestamp 1663859327
transform 1 0 96768 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1850
timestamp 1663859327
transform 1 0 104720 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1851
timestamp 1663859327
transform 1 0 112672 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1852
timestamp 1663859327
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1853
timestamp 1663859327
transform 1 0 13216 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1854
timestamp 1663859327
transform 1 0 21168 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1855
timestamp 1663859327
transform 1 0 29120 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1856
timestamp 1663859327
transform 1 0 37072 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1857
timestamp 1663859327
transform 1 0 45024 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1858
timestamp 1663859327
transform 1 0 52976 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1859
timestamp 1663859327
transform 1 0 60928 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1860
timestamp 1663859327
transform 1 0 68880 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1861
timestamp 1663859327
transform 1 0 76832 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1862
timestamp 1663859327
transform 1 0 84784 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1863
timestamp 1663859327
transform 1 0 92736 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1864
timestamp 1663859327
transform 1 0 100688 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1865
timestamp 1663859327
transform 1 0 108640 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1866
timestamp 1663859327
transform 1 0 116592 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1867
timestamp 1663859327
transform 1 0 9296 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1868
timestamp 1663859327
transform 1 0 17248 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1869
timestamp 1663859327
transform 1 0 25200 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1870
timestamp 1663859327
transform 1 0 33152 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1871
timestamp 1663859327
transform 1 0 41104 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1872
timestamp 1663859327
transform 1 0 49056 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1873
timestamp 1663859327
transform 1 0 57008 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1874
timestamp 1663859327
transform 1 0 64960 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1875
timestamp 1663859327
transform 1 0 72912 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1876
timestamp 1663859327
transform 1 0 80864 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1877
timestamp 1663859327
transform 1 0 88816 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1878
timestamp 1663859327
transform 1 0 96768 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1879
timestamp 1663859327
transform 1 0 104720 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1880
timestamp 1663859327
transform 1 0 112672 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1881
timestamp 1663859327
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1882
timestamp 1663859327
transform 1 0 13216 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1883
timestamp 1663859327
transform 1 0 21168 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1884
timestamp 1663859327
transform 1 0 29120 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1885
timestamp 1663859327
transform 1 0 37072 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1886
timestamp 1663859327
transform 1 0 45024 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1887
timestamp 1663859327
transform 1 0 52976 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1888
timestamp 1663859327
transform 1 0 60928 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1889
timestamp 1663859327
transform 1 0 68880 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1890
timestamp 1663859327
transform 1 0 76832 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1891
timestamp 1663859327
transform 1 0 84784 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1892
timestamp 1663859327
transform 1 0 92736 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1893
timestamp 1663859327
transform 1 0 100688 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1894
timestamp 1663859327
transform 1 0 108640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1895
timestamp 1663859327
transform 1 0 116592 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1896
timestamp 1663859327
transform 1 0 9296 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1897
timestamp 1663859327
transform 1 0 17248 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1898
timestamp 1663859327
transform 1 0 25200 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1899
timestamp 1663859327
transform 1 0 33152 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1900
timestamp 1663859327
transform 1 0 41104 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1901
timestamp 1663859327
transform 1 0 49056 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1902
timestamp 1663859327
transform 1 0 57008 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1903
timestamp 1663859327
transform 1 0 64960 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1904
timestamp 1663859327
transform 1 0 72912 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1905
timestamp 1663859327
transform 1 0 80864 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1906
timestamp 1663859327
transform 1 0 88816 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1907
timestamp 1663859327
transform 1 0 96768 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1908
timestamp 1663859327
transform 1 0 104720 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1909
timestamp 1663859327
transform 1 0 112672 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1910
timestamp 1663859327
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1911
timestamp 1663859327
transform 1 0 13216 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1912
timestamp 1663859327
transform 1 0 21168 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1913
timestamp 1663859327
transform 1 0 29120 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1914
timestamp 1663859327
transform 1 0 37072 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1915
timestamp 1663859327
transform 1 0 45024 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1916
timestamp 1663859327
transform 1 0 52976 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1917
timestamp 1663859327
transform 1 0 60928 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1918
timestamp 1663859327
transform 1 0 68880 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1919
timestamp 1663859327
transform 1 0 76832 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1920
timestamp 1663859327
transform 1 0 84784 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1921
timestamp 1663859327
transform 1 0 92736 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1922
timestamp 1663859327
transform 1 0 100688 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1923
timestamp 1663859327
transform 1 0 108640 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1924
timestamp 1663859327
transform 1 0 116592 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1925
timestamp 1663859327
transform 1 0 9296 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1926
timestamp 1663859327
transform 1 0 17248 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1927
timestamp 1663859327
transform 1 0 25200 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1928
timestamp 1663859327
transform 1 0 33152 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1929
timestamp 1663859327
transform 1 0 41104 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1930
timestamp 1663859327
transform 1 0 49056 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1931
timestamp 1663859327
transform 1 0 57008 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1932
timestamp 1663859327
transform 1 0 64960 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1933
timestamp 1663859327
transform 1 0 72912 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1934
timestamp 1663859327
transform 1 0 80864 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1935
timestamp 1663859327
transform 1 0 88816 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1936
timestamp 1663859327
transform 1 0 96768 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1937
timestamp 1663859327
transform 1 0 104720 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1938
timestamp 1663859327
transform 1 0 112672 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1939
timestamp 1663859327
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1940
timestamp 1663859327
transform 1 0 13216 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1941
timestamp 1663859327
transform 1 0 21168 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1942
timestamp 1663859327
transform 1 0 29120 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1943
timestamp 1663859327
transform 1 0 37072 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1944
timestamp 1663859327
transform 1 0 45024 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1945
timestamp 1663859327
transform 1 0 52976 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1946
timestamp 1663859327
transform 1 0 60928 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1947
timestamp 1663859327
transform 1 0 68880 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1948
timestamp 1663859327
transform 1 0 76832 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1949
timestamp 1663859327
transform 1 0 84784 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1950
timestamp 1663859327
transform 1 0 92736 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1951
timestamp 1663859327
transform 1 0 100688 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1952
timestamp 1663859327
transform 1 0 108640 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1953
timestamp 1663859327
transform 1 0 116592 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1954
timestamp 1663859327
transform 1 0 9296 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1955
timestamp 1663859327
transform 1 0 17248 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1956
timestamp 1663859327
transform 1 0 25200 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1957
timestamp 1663859327
transform 1 0 33152 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1958
timestamp 1663859327
transform 1 0 41104 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1959
timestamp 1663859327
transform 1 0 49056 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1960
timestamp 1663859327
transform 1 0 57008 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1961
timestamp 1663859327
transform 1 0 64960 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1962
timestamp 1663859327
transform 1 0 72912 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1963
timestamp 1663859327
transform 1 0 80864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1964
timestamp 1663859327
transform 1 0 88816 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1965
timestamp 1663859327
transform 1 0 96768 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1966
timestamp 1663859327
transform 1 0 104720 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1967
timestamp 1663859327
transform 1 0 112672 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1968
timestamp 1663859327
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1969
timestamp 1663859327
transform 1 0 13216 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1970
timestamp 1663859327
transform 1 0 21168 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1971
timestamp 1663859327
transform 1 0 29120 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1972
timestamp 1663859327
transform 1 0 37072 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1973
timestamp 1663859327
transform 1 0 45024 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1974
timestamp 1663859327
transform 1 0 52976 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1975
timestamp 1663859327
transform 1 0 60928 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1976
timestamp 1663859327
transform 1 0 68880 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1977
timestamp 1663859327
transform 1 0 76832 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1978
timestamp 1663859327
transform 1 0 84784 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1979
timestamp 1663859327
transform 1 0 92736 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1980
timestamp 1663859327
transform 1 0 100688 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1981
timestamp 1663859327
transform 1 0 108640 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1982
timestamp 1663859327
transform 1 0 116592 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1983
timestamp 1663859327
transform 1 0 9296 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1984
timestamp 1663859327
transform 1 0 17248 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1985
timestamp 1663859327
transform 1 0 25200 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1986
timestamp 1663859327
transform 1 0 33152 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1987
timestamp 1663859327
transform 1 0 41104 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1988
timestamp 1663859327
transform 1 0 49056 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1989
timestamp 1663859327
transform 1 0 57008 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1990
timestamp 1663859327
transform 1 0 64960 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1991
timestamp 1663859327
transform 1 0 72912 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1992
timestamp 1663859327
transform 1 0 80864 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1993
timestamp 1663859327
transform 1 0 88816 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1994
timestamp 1663859327
transform 1 0 96768 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1995
timestamp 1663859327
transform 1 0 104720 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1996
timestamp 1663859327
transform 1 0 112672 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1997
timestamp 1663859327
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1998
timestamp 1663859327
transform 1 0 13216 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1999
timestamp 1663859327
transform 1 0 21168 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2000
timestamp 1663859327
transform 1 0 29120 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2001
timestamp 1663859327
transform 1 0 37072 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2002
timestamp 1663859327
transform 1 0 45024 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2003
timestamp 1663859327
transform 1 0 52976 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2004
timestamp 1663859327
transform 1 0 60928 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2005
timestamp 1663859327
transform 1 0 68880 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2006
timestamp 1663859327
transform 1 0 76832 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2007
timestamp 1663859327
transform 1 0 84784 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2008
timestamp 1663859327
transform 1 0 92736 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2009
timestamp 1663859327
transform 1 0 100688 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2010
timestamp 1663859327
transform 1 0 108640 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2011
timestamp 1663859327
transform 1 0 116592 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2012
timestamp 1663859327
transform 1 0 9296 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2013
timestamp 1663859327
transform 1 0 17248 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2014
timestamp 1663859327
transform 1 0 25200 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2015
timestamp 1663859327
transform 1 0 33152 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2016
timestamp 1663859327
transform 1 0 41104 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2017
timestamp 1663859327
transform 1 0 49056 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2018
timestamp 1663859327
transform 1 0 57008 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2019
timestamp 1663859327
transform 1 0 64960 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2020
timestamp 1663859327
transform 1 0 72912 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2021
timestamp 1663859327
transform 1 0 80864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2022
timestamp 1663859327
transform 1 0 88816 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2023
timestamp 1663859327
transform 1 0 96768 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2024
timestamp 1663859327
transform 1 0 104720 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2025
timestamp 1663859327
transform 1 0 112672 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2026
timestamp 1663859327
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2027
timestamp 1663859327
transform 1 0 13216 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2028
timestamp 1663859327
transform 1 0 21168 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2029
timestamp 1663859327
transform 1 0 29120 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2030
timestamp 1663859327
transform 1 0 37072 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2031
timestamp 1663859327
transform 1 0 45024 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2032
timestamp 1663859327
transform 1 0 52976 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2033
timestamp 1663859327
transform 1 0 60928 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2034
timestamp 1663859327
transform 1 0 68880 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2035
timestamp 1663859327
transform 1 0 76832 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2036
timestamp 1663859327
transform 1 0 84784 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2037
timestamp 1663859327
transform 1 0 92736 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2038
timestamp 1663859327
transform 1 0 100688 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2039
timestamp 1663859327
transform 1 0 108640 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2040
timestamp 1663859327
transform 1 0 116592 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2041
timestamp 1663859327
transform 1 0 9296 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2042
timestamp 1663859327
transform 1 0 17248 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2043
timestamp 1663859327
transform 1 0 25200 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2044
timestamp 1663859327
transform 1 0 33152 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2045
timestamp 1663859327
transform 1 0 41104 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2046
timestamp 1663859327
transform 1 0 49056 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2047
timestamp 1663859327
transform 1 0 57008 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2048
timestamp 1663859327
transform 1 0 64960 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2049
timestamp 1663859327
transform 1 0 72912 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2050
timestamp 1663859327
transform 1 0 80864 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2051
timestamp 1663859327
transform 1 0 88816 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2052
timestamp 1663859327
transform 1 0 96768 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2053
timestamp 1663859327
transform 1 0 104720 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2054
timestamp 1663859327
transform 1 0 112672 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2055
timestamp 1663859327
transform 1 0 5264 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2056
timestamp 1663859327
transform 1 0 13216 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2057
timestamp 1663859327
transform 1 0 21168 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2058
timestamp 1663859327
transform 1 0 29120 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2059
timestamp 1663859327
transform 1 0 37072 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2060
timestamp 1663859327
transform 1 0 45024 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2061
timestamp 1663859327
transform 1 0 52976 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2062
timestamp 1663859327
transform 1 0 60928 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2063
timestamp 1663859327
transform 1 0 68880 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2064
timestamp 1663859327
transform 1 0 76832 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2065
timestamp 1663859327
transform 1 0 84784 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2066
timestamp 1663859327
transform 1 0 92736 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2067
timestamp 1663859327
transform 1 0 100688 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2068
timestamp 1663859327
transform 1 0 108640 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2069
timestamp 1663859327
transform 1 0 116592 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2070
timestamp 1663859327
transform 1 0 9296 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2071
timestamp 1663859327
transform 1 0 17248 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2072
timestamp 1663859327
transform 1 0 25200 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2073
timestamp 1663859327
transform 1 0 33152 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2074
timestamp 1663859327
transform 1 0 41104 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2075
timestamp 1663859327
transform 1 0 49056 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2076
timestamp 1663859327
transform 1 0 57008 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2077
timestamp 1663859327
transform 1 0 64960 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2078
timestamp 1663859327
transform 1 0 72912 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2079
timestamp 1663859327
transform 1 0 80864 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2080
timestamp 1663859327
transform 1 0 88816 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2081
timestamp 1663859327
transform 1 0 96768 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2082
timestamp 1663859327
transform 1 0 104720 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2083
timestamp 1663859327
transform 1 0 112672 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2084
timestamp 1663859327
transform 1 0 5264 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2085
timestamp 1663859327
transform 1 0 13216 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2086
timestamp 1663859327
transform 1 0 21168 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2087
timestamp 1663859327
transform 1 0 29120 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2088
timestamp 1663859327
transform 1 0 37072 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2089
timestamp 1663859327
transform 1 0 45024 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2090
timestamp 1663859327
transform 1 0 52976 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2091
timestamp 1663859327
transform 1 0 60928 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2092
timestamp 1663859327
transform 1 0 68880 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2093
timestamp 1663859327
transform 1 0 76832 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2094
timestamp 1663859327
transform 1 0 84784 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2095
timestamp 1663859327
transform 1 0 92736 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2096
timestamp 1663859327
transform 1 0 100688 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2097
timestamp 1663859327
transform 1 0 108640 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2098
timestamp 1663859327
transform 1 0 116592 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2099
timestamp 1663859327
transform 1 0 9296 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2100
timestamp 1663859327
transform 1 0 17248 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2101
timestamp 1663859327
transform 1 0 25200 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2102
timestamp 1663859327
transform 1 0 33152 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2103
timestamp 1663859327
transform 1 0 41104 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2104
timestamp 1663859327
transform 1 0 49056 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2105
timestamp 1663859327
transform 1 0 57008 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2106
timestamp 1663859327
transform 1 0 64960 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2107
timestamp 1663859327
transform 1 0 72912 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2108
timestamp 1663859327
transform 1 0 80864 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2109
timestamp 1663859327
transform 1 0 88816 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2110
timestamp 1663859327
transform 1 0 96768 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2111
timestamp 1663859327
transform 1 0 104720 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2112
timestamp 1663859327
transform 1 0 112672 0 -1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2113
timestamp 1663859327
transform 1 0 5264 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2114
timestamp 1663859327
transform 1 0 13216 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2115
timestamp 1663859327
transform 1 0 21168 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2116
timestamp 1663859327
transform 1 0 29120 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2117
timestamp 1663859327
transform 1 0 37072 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2118
timestamp 1663859327
transform 1 0 45024 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2119
timestamp 1663859327
transform 1 0 52976 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2120
timestamp 1663859327
transform 1 0 60928 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2121
timestamp 1663859327
transform 1 0 68880 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2122
timestamp 1663859327
transform 1 0 76832 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2123
timestamp 1663859327
transform 1 0 84784 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2124
timestamp 1663859327
transform 1 0 92736 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2125
timestamp 1663859327
transform 1 0 100688 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2126
timestamp 1663859327
transform 1 0 108640 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2127
timestamp 1663859327
transform 1 0 116592 0 1 98784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2128
timestamp 1663859327
transform 1 0 9296 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2129
timestamp 1663859327
transform 1 0 17248 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2130
timestamp 1663859327
transform 1 0 25200 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2131
timestamp 1663859327
transform 1 0 33152 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2132
timestamp 1663859327
transform 1 0 41104 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2133
timestamp 1663859327
transform 1 0 49056 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2134
timestamp 1663859327
transform 1 0 57008 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2135
timestamp 1663859327
transform 1 0 64960 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2136
timestamp 1663859327
transform 1 0 72912 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2137
timestamp 1663859327
transform 1 0 80864 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2138
timestamp 1663859327
transform 1 0 88816 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2139
timestamp 1663859327
transform 1 0 96768 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2140
timestamp 1663859327
transform 1 0 104720 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2141
timestamp 1663859327
transform 1 0 112672 0 -1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2142
timestamp 1663859327
transform 1 0 5264 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2143
timestamp 1663859327
transform 1 0 13216 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2144
timestamp 1663859327
transform 1 0 21168 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2145
timestamp 1663859327
transform 1 0 29120 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2146
timestamp 1663859327
transform 1 0 37072 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2147
timestamp 1663859327
transform 1 0 45024 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2148
timestamp 1663859327
transform 1 0 52976 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2149
timestamp 1663859327
transform 1 0 60928 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2150
timestamp 1663859327
transform 1 0 68880 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2151
timestamp 1663859327
transform 1 0 76832 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2152
timestamp 1663859327
transform 1 0 84784 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2153
timestamp 1663859327
transform 1 0 92736 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2154
timestamp 1663859327
transform 1 0 100688 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2155
timestamp 1663859327
transform 1 0 108640 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2156
timestamp 1663859327
transform 1 0 116592 0 1 100352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2157
timestamp 1663859327
transform 1 0 9296 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2158
timestamp 1663859327
transform 1 0 17248 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2159
timestamp 1663859327
transform 1 0 25200 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2160
timestamp 1663859327
transform 1 0 33152 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2161
timestamp 1663859327
transform 1 0 41104 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2162
timestamp 1663859327
transform 1 0 49056 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2163
timestamp 1663859327
transform 1 0 57008 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2164
timestamp 1663859327
transform 1 0 64960 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2165
timestamp 1663859327
transform 1 0 72912 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2166
timestamp 1663859327
transform 1 0 80864 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2167
timestamp 1663859327
transform 1 0 88816 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2168
timestamp 1663859327
transform 1 0 96768 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2169
timestamp 1663859327
transform 1 0 104720 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2170
timestamp 1663859327
transform 1 0 112672 0 -1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2171
timestamp 1663859327
transform 1 0 5264 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2172
timestamp 1663859327
transform 1 0 13216 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2173
timestamp 1663859327
transform 1 0 21168 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2174
timestamp 1663859327
transform 1 0 29120 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2175
timestamp 1663859327
transform 1 0 37072 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2176
timestamp 1663859327
transform 1 0 45024 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2177
timestamp 1663859327
transform 1 0 52976 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2178
timestamp 1663859327
transform 1 0 60928 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2179
timestamp 1663859327
transform 1 0 68880 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2180
timestamp 1663859327
transform 1 0 76832 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2181
timestamp 1663859327
transform 1 0 84784 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2182
timestamp 1663859327
transform 1 0 92736 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2183
timestamp 1663859327
transform 1 0 100688 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2184
timestamp 1663859327
transform 1 0 108640 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2185
timestamp 1663859327
transform 1 0 116592 0 1 101920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2186
timestamp 1663859327
transform 1 0 9296 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2187
timestamp 1663859327
transform 1 0 17248 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2188
timestamp 1663859327
transform 1 0 25200 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2189
timestamp 1663859327
transform 1 0 33152 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2190
timestamp 1663859327
transform 1 0 41104 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2191
timestamp 1663859327
transform 1 0 49056 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2192
timestamp 1663859327
transform 1 0 57008 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2193
timestamp 1663859327
transform 1 0 64960 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2194
timestamp 1663859327
transform 1 0 72912 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2195
timestamp 1663859327
transform 1 0 80864 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2196
timestamp 1663859327
transform 1 0 88816 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2197
timestamp 1663859327
transform 1 0 96768 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2198
timestamp 1663859327
transform 1 0 104720 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2199
timestamp 1663859327
transform 1 0 112672 0 -1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2200
timestamp 1663859327
transform 1 0 5264 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2201
timestamp 1663859327
transform 1 0 13216 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2202
timestamp 1663859327
transform 1 0 21168 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2203
timestamp 1663859327
transform 1 0 29120 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2204
timestamp 1663859327
transform 1 0 37072 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2205
timestamp 1663859327
transform 1 0 45024 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2206
timestamp 1663859327
transform 1 0 52976 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2207
timestamp 1663859327
transform 1 0 60928 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2208
timestamp 1663859327
transform 1 0 68880 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2209
timestamp 1663859327
transform 1 0 76832 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2210
timestamp 1663859327
transform 1 0 84784 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2211
timestamp 1663859327
transform 1 0 92736 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2212
timestamp 1663859327
transform 1 0 100688 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2213
timestamp 1663859327
transform 1 0 108640 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2214
timestamp 1663859327
transform 1 0 116592 0 1 103488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2215
timestamp 1663859327
transform 1 0 9296 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2216
timestamp 1663859327
transform 1 0 17248 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2217
timestamp 1663859327
transform 1 0 25200 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2218
timestamp 1663859327
transform 1 0 33152 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2219
timestamp 1663859327
transform 1 0 41104 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2220
timestamp 1663859327
transform 1 0 49056 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2221
timestamp 1663859327
transform 1 0 57008 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2222
timestamp 1663859327
transform 1 0 64960 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2223
timestamp 1663859327
transform 1 0 72912 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2224
timestamp 1663859327
transform 1 0 80864 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2225
timestamp 1663859327
transform 1 0 88816 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2226
timestamp 1663859327
transform 1 0 96768 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2227
timestamp 1663859327
transform 1 0 104720 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2228
timestamp 1663859327
transform 1 0 112672 0 -1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2229
timestamp 1663859327
transform 1 0 5264 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2230
timestamp 1663859327
transform 1 0 13216 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2231
timestamp 1663859327
transform 1 0 21168 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2232
timestamp 1663859327
transform 1 0 29120 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2233
timestamp 1663859327
transform 1 0 37072 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2234
timestamp 1663859327
transform 1 0 45024 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2235
timestamp 1663859327
transform 1 0 52976 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2236
timestamp 1663859327
transform 1 0 60928 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2237
timestamp 1663859327
transform 1 0 68880 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2238
timestamp 1663859327
transform 1 0 76832 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2239
timestamp 1663859327
transform 1 0 84784 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2240
timestamp 1663859327
transform 1 0 92736 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2241
timestamp 1663859327
transform 1 0 100688 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2242
timestamp 1663859327
transform 1 0 108640 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2243
timestamp 1663859327
transform 1 0 116592 0 1 105056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2244
timestamp 1663859327
transform 1 0 9296 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2245
timestamp 1663859327
transform 1 0 17248 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2246
timestamp 1663859327
transform 1 0 25200 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2247
timestamp 1663859327
transform 1 0 33152 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2248
timestamp 1663859327
transform 1 0 41104 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2249
timestamp 1663859327
transform 1 0 49056 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2250
timestamp 1663859327
transform 1 0 57008 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2251
timestamp 1663859327
transform 1 0 64960 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2252
timestamp 1663859327
transform 1 0 72912 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2253
timestamp 1663859327
transform 1 0 80864 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2254
timestamp 1663859327
transform 1 0 88816 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2255
timestamp 1663859327
transform 1 0 96768 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2256
timestamp 1663859327
transform 1 0 104720 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2257
timestamp 1663859327
transform 1 0 112672 0 -1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2258
timestamp 1663859327
transform 1 0 5264 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2259
timestamp 1663859327
transform 1 0 13216 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2260
timestamp 1663859327
transform 1 0 21168 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2261
timestamp 1663859327
transform 1 0 29120 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2262
timestamp 1663859327
transform 1 0 37072 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2263
timestamp 1663859327
transform 1 0 45024 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2264
timestamp 1663859327
transform 1 0 52976 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2265
timestamp 1663859327
transform 1 0 60928 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2266
timestamp 1663859327
transform 1 0 68880 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2267
timestamp 1663859327
transform 1 0 76832 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2268
timestamp 1663859327
transform 1 0 84784 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2269
timestamp 1663859327
transform 1 0 92736 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2270
timestamp 1663859327
transform 1 0 100688 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2271
timestamp 1663859327
transform 1 0 108640 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2272
timestamp 1663859327
transform 1 0 116592 0 1 106624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2273
timestamp 1663859327
transform 1 0 9296 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2274
timestamp 1663859327
transform 1 0 17248 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2275
timestamp 1663859327
transform 1 0 25200 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2276
timestamp 1663859327
transform 1 0 33152 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2277
timestamp 1663859327
transform 1 0 41104 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2278
timestamp 1663859327
transform 1 0 49056 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2279
timestamp 1663859327
transform 1 0 57008 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2280
timestamp 1663859327
transform 1 0 64960 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2281
timestamp 1663859327
transform 1 0 72912 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2282
timestamp 1663859327
transform 1 0 80864 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2283
timestamp 1663859327
transform 1 0 88816 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2284
timestamp 1663859327
transform 1 0 96768 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2285
timestamp 1663859327
transform 1 0 104720 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2286
timestamp 1663859327
transform 1 0 112672 0 -1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2287
timestamp 1663859327
transform 1 0 5264 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2288
timestamp 1663859327
transform 1 0 13216 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2289
timestamp 1663859327
transform 1 0 21168 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2290
timestamp 1663859327
transform 1 0 29120 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2291
timestamp 1663859327
transform 1 0 37072 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2292
timestamp 1663859327
transform 1 0 45024 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2293
timestamp 1663859327
transform 1 0 52976 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2294
timestamp 1663859327
transform 1 0 60928 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2295
timestamp 1663859327
transform 1 0 68880 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2296
timestamp 1663859327
transform 1 0 76832 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2297
timestamp 1663859327
transform 1 0 84784 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2298
timestamp 1663859327
transform 1 0 92736 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2299
timestamp 1663859327
transform 1 0 100688 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2300
timestamp 1663859327
transform 1 0 108640 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2301
timestamp 1663859327
transform 1 0 116592 0 1 108192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2302
timestamp 1663859327
transform 1 0 9296 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2303
timestamp 1663859327
transform 1 0 17248 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2304
timestamp 1663859327
transform 1 0 25200 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2305
timestamp 1663859327
transform 1 0 33152 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2306
timestamp 1663859327
transform 1 0 41104 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2307
timestamp 1663859327
transform 1 0 49056 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2308
timestamp 1663859327
transform 1 0 57008 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2309
timestamp 1663859327
transform 1 0 64960 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2310
timestamp 1663859327
transform 1 0 72912 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2311
timestamp 1663859327
transform 1 0 80864 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2312
timestamp 1663859327
transform 1 0 88816 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2313
timestamp 1663859327
transform 1 0 96768 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2314
timestamp 1663859327
transform 1 0 104720 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2315
timestamp 1663859327
transform 1 0 112672 0 -1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2316
timestamp 1663859327
transform 1 0 5264 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2317
timestamp 1663859327
transform 1 0 13216 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2318
timestamp 1663859327
transform 1 0 21168 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2319
timestamp 1663859327
transform 1 0 29120 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2320
timestamp 1663859327
transform 1 0 37072 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2321
timestamp 1663859327
transform 1 0 45024 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2322
timestamp 1663859327
transform 1 0 52976 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2323
timestamp 1663859327
transform 1 0 60928 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2324
timestamp 1663859327
transform 1 0 68880 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2325
timestamp 1663859327
transform 1 0 76832 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2326
timestamp 1663859327
transform 1 0 84784 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2327
timestamp 1663859327
transform 1 0 92736 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2328
timestamp 1663859327
transform 1 0 100688 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2329
timestamp 1663859327
transform 1 0 108640 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2330
timestamp 1663859327
transform 1 0 116592 0 1 109760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2331
timestamp 1663859327
transform 1 0 9296 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2332
timestamp 1663859327
transform 1 0 17248 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2333
timestamp 1663859327
transform 1 0 25200 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2334
timestamp 1663859327
transform 1 0 33152 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2335
timestamp 1663859327
transform 1 0 41104 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2336
timestamp 1663859327
transform 1 0 49056 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2337
timestamp 1663859327
transform 1 0 57008 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2338
timestamp 1663859327
transform 1 0 64960 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2339
timestamp 1663859327
transform 1 0 72912 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2340
timestamp 1663859327
transform 1 0 80864 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2341
timestamp 1663859327
transform 1 0 88816 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2342
timestamp 1663859327
transform 1 0 96768 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2343
timestamp 1663859327
transform 1 0 104720 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2344
timestamp 1663859327
transform 1 0 112672 0 -1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2345
timestamp 1663859327
transform 1 0 5264 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2346
timestamp 1663859327
transform 1 0 13216 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2347
timestamp 1663859327
transform 1 0 21168 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2348
timestamp 1663859327
transform 1 0 29120 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2349
timestamp 1663859327
transform 1 0 37072 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2350
timestamp 1663859327
transform 1 0 45024 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2351
timestamp 1663859327
transform 1 0 52976 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2352
timestamp 1663859327
transform 1 0 60928 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2353
timestamp 1663859327
transform 1 0 68880 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2354
timestamp 1663859327
transform 1 0 76832 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2355
timestamp 1663859327
transform 1 0 84784 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2356
timestamp 1663859327
transform 1 0 92736 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2357
timestamp 1663859327
transform 1 0 100688 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2358
timestamp 1663859327
transform 1 0 108640 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2359
timestamp 1663859327
transform 1 0 116592 0 1 111328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2360
timestamp 1663859327
transform 1 0 9296 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2361
timestamp 1663859327
transform 1 0 17248 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2362
timestamp 1663859327
transform 1 0 25200 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2363
timestamp 1663859327
transform 1 0 33152 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2364
timestamp 1663859327
transform 1 0 41104 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2365
timestamp 1663859327
transform 1 0 49056 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2366
timestamp 1663859327
transform 1 0 57008 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2367
timestamp 1663859327
transform 1 0 64960 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2368
timestamp 1663859327
transform 1 0 72912 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2369
timestamp 1663859327
transform 1 0 80864 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2370
timestamp 1663859327
transform 1 0 88816 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2371
timestamp 1663859327
transform 1 0 96768 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2372
timestamp 1663859327
transform 1 0 104720 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2373
timestamp 1663859327
transform 1 0 112672 0 -1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2374
timestamp 1663859327
transform 1 0 5264 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2375
timestamp 1663859327
transform 1 0 13216 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2376
timestamp 1663859327
transform 1 0 21168 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2377
timestamp 1663859327
transform 1 0 29120 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2378
timestamp 1663859327
transform 1 0 37072 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2379
timestamp 1663859327
transform 1 0 45024 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2380
timestamp 1663859327
transform 1 0 52976 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2381
timestamp 1663859327
transform 1 0 60928 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2382
timestamp 1663859327
transform 1 0 68880 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2383
timestamp 1663859327
transform 1 0 76832 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2384
timestamp 1663859327
transform 1 0 84784 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2385
timestamp 1663859327
transform 1 0 92736 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2386
timestamp 1663859327
transform 1 0 100688 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2387
timestamp 1663859327
transform 1 0 108640 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2388
timestamp 1663859327
transform 1 0 116592 0 1 112896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2389
timestamp 1663859327
transform 1 0 9296 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2390
timestamp 1663859327
transform 1 0 17248 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2391
timestamp 1663859327
transform 1 0 25200 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2392
timestamp 1663859327
transform 1 0 33152 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2393
timestamp 1663859327
transform 1 0 41104 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2394
timestamp 1663859327
transform 1 0 49056 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2395
timestamp 1663859327
transform 1 0 57008 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2396
timestamp 1663859327
transform 1 0 64960 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2397
timestamp 1663859327
transform 1 0 72912 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2398
timestamp 1663859327
transform 1 0 80864 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2399
timestamp 1663859327
transform 1 0 88816 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2400
timestamp 1663859327
transform 1 0 96768 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2401
timestamp 1663859327
transform 1 0 104720 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2402
timestamp 1663859327
transform 1 0 112672 0 -1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2403
timestamp 1663859327
transform 1 0 5264 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2404
timestamp 1663859327
transform 1 0 13216 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2405
timestamp 1663859327
transform 1 0 21168 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2406
timestamp 1663859327
transform 1 0 29120 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2407
timestamp 1663859327
transform 1 0 37072 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2408
timestamp 1663859327
transform 1 0 45024 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2409
timestamp 1663859327
transform 1 0 52976 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2410
timestamp 1663859327
transform 1 0 60928 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2411
timestamp 1663859327
transform 1 0 68880 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2412
timestamp 1663859327
transform 1 0 76832 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2413
timestamp 1663859327
transform 1 0 84784 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2414
timestamp 1663859327
transform 1 0 92736 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2415
timestamp 1663859327
transform 1 0 100688 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2416
timestamp 1663859327
transform 1 0 108640 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2417
timestamp 1663859327
transform 1 0 116592 0 1 114464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2418
timestamp 1663859327
transform 1 0 9296 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2419
timestamp 1663859327
transform 1 0 17248 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2420
timestamp 1663859327
transform 1 0 25200 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2421
timestamp 1663859327
transform 1 0 33152 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2422
timestamp 1663859327
transform 1 0 41104 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2423
timestamp 1663859327
transform 1 0 49056 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2424
timestamp 1663859327
transform 1 0 57008 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2425
timestamp 1663859327
transform 1 0 64960 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2426
timestamp 1663859327
transform 1 0 72912 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2427
timestamp 1663859327
transform 1 0 80864 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2428
timestamp 1663859327
transform 1 0 88816 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2429
timestamp 1663859327
transform 1 0 96768 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2430
timestamp 1663859327
transform 1 0 104720 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2431
timestamp 1663859327
transform 1 0 112672 0 -1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2432
timestamp 1663859327
transform 1 0 5264 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2433
timestamp 1663859327
transform 1 0 13216 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2434
timestamp 1663859327
transform 1 0 21168 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2435
timestamp 1663859327
transform 1 0 29120 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2436
timestamp 1663859327
transform 1 0 37072 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2437
timestamp 1663859327
transform 1 0 45024 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2438
timestamp 1663859327
transform 1 0 52976 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2439
timestamp 1663859327
transform 1 0 60928 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2440
timestamp 1663859327
transform 1 0 68880 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2441
timestamp 1663859327
transform 1 0 76832 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2442
timestamp 1663859327
transform 1 0 84784 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2443
timestamp 1663859327
transform 1 0 92736 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2444
timestamp 1663859327
transform 1 0 100688 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2445
timestamp 1663859327
transform 1 0 108640 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2446
timestamp 1663859327
transform 1 0 116592 0 1 116032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2447
timestamp 1663859327
transform 1 0 9296 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2448
timestamp 1663859327
transform 1 0 17248 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2449
timestamp 1663859327
transform 1 0 25200 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2450
timestamp 1663859327
transform 1 0 33152 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2451
timestamp 1663859327
transform 1 0 41104 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2452
timestamp 1663859327
transform 1 0 49056 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2453
timestamp 1663859327
transform 1 0 57008 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2454
timestamp 1663859327
transform 1 0 64960 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2455
timestamp 1663859327
transform 1 0 72912 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2456
timestamp 1663859327
transform 1 0 80864 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2457
timestamp 1663859327
transform 1 0 88816 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2458
timestamp 1663859327
transform 1 0 96768 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2459
timestamp 1663859327
transform 1 0 104720 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2460
timestamp 1663859327
transform 1 0 112672 0 -1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2461
timestamp 1663859327
transform 1 0 5264 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2462
timestamp 1663859327
transform 1 0 13216 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2463
timestamp 1663859327
transform 1 0 21168 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2464
timestamp 1663859327
transform 1 0 29120 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2465
timestamp 1663859327
transform 1 0 37072 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2466
timestamp 1663859327
transform 1 0 45024 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2467
timestamp 1663859327
transform 1 0 52976 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2468
timestamp 1663859327
transform 1 0 60928 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2469
timestamp 1663859327
transform 1 0 68880 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2470
timestamp 1663859327
transform 1 0 76832 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2471
timestamp 1663859327
transform 1 0 84784 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2472
timestamp 1663859327
transform 1 0 92736 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2473
timestamp 1663859327
transform 1 0 100688 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2474
timestamp 1663859327
transform 1 0 108640 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2475
timestamp 1663859327
transform 1 0 116592 0 1 117600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2476
timestamp 1663859327
transform 1 0 9296 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2477
timestamp 1663859327
transform 1 0 17248 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2478
timestamp 1663859327
transform 1 0 25200 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2479
timestamp 1663859327
transform 1 0 33152 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2480
timestamp 1663859327
transform 1 0 41104 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2481
timestamp 1663859327
transform 1 0 49056 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2482
timestamp 1663859327
transform 1 0 57008 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2483
timestamp 1663859327
transform 1 0 64960 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2484
timestamp 1663859327
transform 1 0 72912 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2485
timestamp 1663859327
transform 1 0 80864 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2486
timestamp 1663859327
transform 1 0 88816 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2487
timestamp 1663859327
transform 1 0 96768 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2488
timestamp 1663859327
transform 1 0 104720 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2489
timestamp 1663859327
transform 1 0 112672 0 -1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2490
timestamp 1663859327
transform 1 0 5264 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2491
timestamp 1663859327
transform 1 0 13216 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2492
timestamp 1663859327
transform 1 0 21168 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2493
timestamp 1663859327
transform 1 0 29120 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2494
timestamp 1663859327
transform 1 0 37072 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2495
timestamp 1663859327
transform 1 0 45024 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2496
timestamp 1663859327
transform 1 0 52976 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2497
timestamp 1663859327
transform 1 0 60928 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2498
timestamp 1663859327
transform 1 0 68880 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2499
timestamp 1663859327
transform 1 0 76832 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2500
timestamp 1663859327
transform 1 0 84784 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2501
timestamp 1663859327
transform 1 0 92736 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2502
timestamp 1663859327
transform 1 0 100688 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2503
timestamp 1663859327
transform 1 0 108640 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2504
timestamp 1663859327
transform 1 0 116592 0 1 119168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2505
timestamp 1663859327
transform 1 0 9296 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2506
timestamp 1663859327
transform 1 0 17248 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2507
timestamp 1663859327
transform 1 0 25200 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2508
timestamp 1663859327
transform 1 0 33152 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2509
timestamp 1663859327
transform 1 0 41104 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2510
timestamp 1663859327
transform 1 0 49056 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2511
timestamp 1663859327
transform 1 0 57008 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2512
timestamp 1663859327
transform 1 0 64960 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2513
timestamp 1663859327
transform 1 0 72912 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2514
timestamp 1663859327
transform 1 0 80864 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2515
timestamp 1663859327
transform 1 0 88816 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2516
timestamp 1663859327
transform 1 0 96768 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2517
timestamp 1663859327
transform 1 0 104720 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2518
timestamp 1663859327
transform 1 0 112672 0 -1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2519
timestamp 1663859327
transform 1 0 5264 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2520
timestamp 1663859327
transform 1 0 13216 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2521
timestamp 1663859327
transform 1 0 21168 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2522
timestamp 1663859327
transform 1 0 29120 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2523
timestamp 1663859327
transform 1 0 37072 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2524
timestamp 1663859327
transform 1 0 45024 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2525
timestamp 1663859327
transform 1 0 52976 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2526
timestamp 1663859327
transform 1 0 60928 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2527
timestamp 1663859327
transform 1 0 68880 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2528
timestamp 1663859327
transform 1 0 76832 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2529
timestamp 1663859327
transform 1 0 84784 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2530
timestamp 1663859327
transform 1 0 92736 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2531
timestamp 1663859327
transform 1 0 100688 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2532
timestamp 1663859327
transform 1 0 108640 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2533
timestamp 1663859327
transform 1 0 116592 0 1 120736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2534
timestamp 1663859327
transform 1 0 9296 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2535
timestamp 1663859327
transform 1 0 17248 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2536
timestamp 1663859327
transform 1 0 25200 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2537
timestamp 1663859327
transform 1 0 33152 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2538
timestamp 1663859327
transform 1 0 41104 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2539
timestamp 1663859327
transform 1 0 49056 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2540
timestamp 1663859327
transform 1 0 57008 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2541
timestamp 1663859327
transform 1 0 64960 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2542
timestamp 1663859327
transform 1 0 72912 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2543
timestamp 1663859327
transform 1 0 80864 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2544
timestamp 1663859327
transform 1 0 88816 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2545
timestamp 1663859327
transform 1 0 96768 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2546
timestamp 1663859327
transform 1 0 104720 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2547
timestamp 1663859327
transform 1 0 112672 0 -1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2548
timestamp 1663859327
transform 1 0 5264 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2549
timestamp 1663859327
transform 1 0 13216 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2550
timestamp 1663859327
transform 1 0 21168 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2551
timestamp 1663859327
transform 1 0 29120 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2552
timestamp 1663859327
transform 1 0 37072 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2553
timestamp 1663859327
transform 1 0 45024 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2554
timestamp 1663859327
transform 1 0 52976 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2555
timestamp 1663859327
transform 1 0 60928 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2556
timestamp 1663859327
transform 1 0 68880 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2557
timestamp 1663859327
transform 1 0 76832 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2558
timestamp 1663859327
transform 1 0 84784 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2559
timestamp 1663859327
transform 1 0 92736 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2560
timestamp 1663859327
transform 1 0 100688 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2561
timestamp 1663859327
transform 1 0 108640 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2562
timestamp 1663859327
transform 1 0 116592 0 1 122304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2563
timestamp 1663859327
transform 1 0 9296 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2564
timestamp 1663859327
transform 1 0 17248 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2565
timestamp 1663859327
transform 1 0 25200 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2566
timestamp 1663859327
transform 1 0 33152 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2567
timestamp 1663859327
transform 1 0 41104 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2568
timestamp 1663859327
transform 1 0 49056 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2569
timestamp 1663859327
transform 1 0 57008 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2570
timestamp 1663859327
transform 1 0 64960 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2571
timestamp 1663859327
transform 1 0 72912 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2572
timestamp 1663859327
transform 1 0 80864 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2573
timestamp 1663859327
transform 1 0 88816 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2574
timestamp 1663859327
transform 1 0 96768 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2575
timestamp 1663859327
transform 1 0 104720 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2576
timestamp 1663859327
transform 1 0 112672 0 -1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2577
timestamp 1663859327
transform 1 0 5264 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2578
timestamp 1663859327
transform 1 0 13216 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2579
timestamp 1663859327
transform 1 0 21168 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2580
timestamp 1663859327
transform 1 0 29120 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2581
timestamp 1663859327
transform 1 0 37072 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2582
timestamp 1663859327
transform 1 0 45024 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2583
timestamp 1663859327
transform 1 0 52976 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2584
timestamp 1663859327
transform 1 0 60928 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2585
timestamp 1663859327
transform 1 0 68880 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2586
timestamp 1663859327
transform 1 0 76832 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2587
timestamp 1663859327
transform 1 0 84784 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2588
timestamp 1663859327
transform 1 0 92736 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2589
timestamp 1663859327
transform 1 0 100688 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2590
timestamp 1663859327
transform 1 0 108640 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2591
timestamp 1663859327
transform 1 0 116592 0 1 123872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2592
timestamp 1663859327
transform 1 0 9296 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2593
timestamp 1663859327
transform 1 0 17248 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2594
timestamp 1663859327
transform 1 0 25200 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2595
timestamp 1663859327
transform 1 0 33152 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2596
timestamp 1663859327
transform 1 0 41104 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2597
timestamp 1663859327
transform 1 0 49056 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2598
timestamp 1663859327
transform 1 0 57008 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2599
timestamp 1663859327
transform 1 0 64960 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2600
timestamp 1663859327
transform 1 0 72912 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2601
timestamp 1663859327
transform 1 0 80864 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2602
timestamp 1663859327
transform 1 0 88816 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2603
timestamp 1663859327
transform 1 0 96768 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2604
timestamp 1663859327
transform 1 0 104720 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2605
timestamp 1663859327
transform 1 0 112672 0 -1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2606
timestamp 1663859327
transform 1 0 5264 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2607
timestamp 1663859327
transform 1 0 13216 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2608
timestamp 1663859327
transform 1 0 21168 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2609
timestamp 1663859327
transform 1 0 29120 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2610
timestamp 1663859327
transform 1 0 37072 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2611
timestamp 1663859327
transform 1 0 45024 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2612
timestamp 1663859327
transform 1 0 52976 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2613
timestamp 1663859327
transform 1 0 60928 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2614
timestamp 1663859327
transform 1 0 68880 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2615
timestamp 1663859327
transform 1 0 76832 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2616
timestamp 1663859327
transform 1 0 84784 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2617
timestamp 1663859327
transform 1 0 92736 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2618
timestamp 1663859327
transform 1 0 100688 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2619
timestamp 1663859327
transform 1 0 108640 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2620
timestamp 1663859327
transform 1 0 116592 0 1 125440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2621
timestamp 1663859327
transform 1 0 9296 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2622
timestamp 1663859327
transform 1 0 17248 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2623
timestamp 1663859327
transform 1 0 25200 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2624
timestamp 1663859327
transform 1 0 33152 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2625
timestamp 1663859327
transform 1 0 41104 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2626
timestamp 1663859327
transform 1 0 49056 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2627
timestamp 1663859327
transform 1 0 57008 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2628
timestamp 1663859327
transform 1 0 64960 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2629
timestamp 1663859327
transform 1 0 72912 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2630
timestamp 1663859327
transform 1 0 80864 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2631
timestamp 1663859327
transform 1 0 88816 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2632
timestamp 1663859327
transform 1 0 96768 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2633
timestamp 1663859327
transform 1 0 104720 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2634
timestamp 1663859327
transform 1 0 112672 0 -1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2635
timestamp 1663859327
transform 1 0 5264 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2636
timestamp 1663859327
transform 1 0 13216 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2637
timestamp 1663859327
transform 1 0 21168 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2638
timestamp 1663859327
transform 1 0 29120 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2639
timestamp 1663859327
transform 1 0 37072 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2640
timestamp 1663859327
transform 1 0 45024 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2641
timestamp 1663859327
transform 1 0 52976 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2642
timestamp 1663859327
transform 1 0 60928 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2643
timestamp 1663859327
transform 1 0 68880 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2644
timestamp 1663859327
transform 1 0 76832 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2645
timestamp 1663859327
transform 1 0 84784 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2646
timestamp 1663859327
transform 1 0 92736 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2647
timestamp 1663859327
transform 1 0 100688 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2648
timestamp 1663859327
transform 1 0 108640 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2649
timestamp 1663859327
transform 1 0 116592 0 1 127008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2650
timestamp 1663859327
transform 1 0 9296 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2651
timestamp 1663859327
transform 1 0 17248 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2652
timestamp 1663859327
transform 1 0 25200 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2653
timestamp 1663859327
transform 1 0 33152 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2654
timestamp 1663859327
transform 1 0 41104 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2655
timestamp 1663859327
transform 1 0 49056 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2656
timestamp 1663859327
transform 1 0 57008 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2657
timestamp 1663859327
transform 1 0 64960 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2658
timestamp 1663859327
transform 1 0 72912 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2659
timestamp 1663859327
transform 1 0 80864 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2660
timestamp 1663859327
transform 1 0 88816 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2661
timestamp 1663859327
transform 1 0 96768 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2662
timestamp 1663859327
transform 1 0 104720 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2663
timestamp 1663859327
transform 1 0 112672 0 -1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2664
timestamp 1663859327
transform 1 0 5264 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2665
timestamp 1663859327
transform 1 0 13216 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2666
timestamp 1663859327
transform 1 0 21168 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2667
timestamp 1663859327
transform 1 0 29120 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2668
timestamp 1663859327
transform 1 0 37072 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2669
timestamp 1663859327
transform 1 0 45024 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2670
timestamp 1663859327
transform 1 0 52976 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2671
timestamp 1663859327
transform 1 0 60928 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2672
timestamp 1663859327
transform 1 0 68880 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2673
timestamp 1663859327
transform 1 0 76832 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2674
timestamp 1663859327
transform 1 0 84784 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2675
timestamp 1663859327
transform 1 0 92736 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2676
timestamp 1663859327
transform 1 0 100688 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2677
timestamp 1663859327
transform 1 0 108640 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2678
timestamp 1663859327
transform 1 0 116592 0 1 128576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2679
timestamp 1663859327
transform 1 0 9296 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2680
timestamp 1663859327
transform 1 0 17248 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2681
timestamp 1663859327
transform 1 0 25200 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2682
timestamp 1663859327
transform 1 0 33152 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2683
timestamp 1663859327
transform 1 0 41104 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2684
timestamp 1663859327
transform 1 0 49056 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2685
timestamp 1663859327
transform 1 0 57008 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2686
timestamp 1663859327
transform 1 0 64960 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2687
timestamp 1663859327
transform 1 0 72912 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2688
timestamp 1663859327
transform 1 0 80864 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2689
timestamp 1663859327
transform 1 0 88816 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2690
timestamp 1663859327
transform 1 0 96768 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2691
timestamp 1663859327
transform 1 0 104720 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2692
timestamp 1663859327
transform 1 0 112672 0 -1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2693
timestamp 1663859327
transform 1 0 5264 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2694
timestamp 1663859327
transform 1 0 13216 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2695
timestamp 1663859327
transform 1 0 21168 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2696
timestamp 1663859327
transform 1 0 29120 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2697
timestamp 1663859327
transform 1 0 37072 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2698
timestamp 1663859327
transform 1 0 45024 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2699
timestamp 1663859327
transform 1 0 52976 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2700
timestamp 1663859327
transform 1 0 60928 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2701
timestamp 1663859327
transform 1 0 68880 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2702
timestamp 1663859327
transform 1 0 76832 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2703
timestamp 1663859327
transform 1 0 84784 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2704
timestamp 1663859327
transform 1 0 92736 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2705
timestamp 1663859327
transform 1 0 100688 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2706
timestamp 1663859327
transform 1 0 108640 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2707
timestamp 1663859327
transform 1 0 116592 0 1 130144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2708
timestamp 1663859327
transform 1 0 9296 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2709
timestamp 1663859327
transform 1 0 17248 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2710
timestamp 1663859327
transform 1 0 25200 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2711
timestamp 1663859327
transform 1 0 33152 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2712
timestamp 1663859327
transform 1 0 41104 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2713
timestamp 1663859327
transform 1 0 49056 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2714
timestamp 1663859327
transform 1 0 57008 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2715
timestamp 1663859327
transform 1 0 64960 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2716
timestamp 1663859327
transform 1 0 72912 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2717
timestamp 1663859327
transform 1 0 80864 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2718
timestamp 1663859327
transform 1 0 88816 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2719
timestamp 1663859327
transform 1 0 96768 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2720
timestamp 1663859327
transform 1 0 104720 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2721
timestamp 1663859327
transform 1 0 112672 0 -1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2722
timestamp 1663859327
transform 1 0 5264 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2723
timestamp 1663859327
transform 1 0 9184 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2724
timestamp 1663859327
transform 1 0 13104 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2725
timestamp 1663859327
transform 1 0 17024 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2726
timestamp 1663859327
transform 1 0 20944 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2727
timestamp 1663859327
transform 1 0 24864 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2728
timestamp 1663859327
transform 1 0 28784 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2729
timestamp 1663859327
transform 1 0 32704 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2730
timestamp 1663859327
transform 1 0 36624 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2731
timestamp 1663859327
transform 1 0 40544 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2732
timestamp 1663859327
transform 1 0 44464 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2733
timestamp 1663859327
transform 1 0 48384 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2734
timestamp 1663859327
transform 1 0 52304 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2735
timestamp 1663859327
transform 1 0 56224 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2736
timestamp 1663859327
transform 1 0 60144 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2737
timestamp 1663859327
transform 1 0 64064 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2738
timestamp 1663859327
transform 1 0 67984 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2739
timestamp 1663859327
transform 1 0 71904 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2740
timestamp 1663859327
transform 1 0 75824 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2741
timestamp 1663859327
transform 1 0 79744 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2742
timestamp 1663859327
transform 1 0 83664 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2743
timestamp 1663859327
transform 1 0 87584 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2744
timestamp 1663859327
transform 1 0 91504 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2745
timestamp 1663859327
transform 1 0 95424 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2746
timestamp 1663859327
transform 1 0 99344 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2747
timestamp 1663859327
transform 1 0 103264 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2748
timestamp 1663859327
transform 1 0 107184 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2749
timestamp 1663859327
transform 1 0 111104 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_2750
timestamp 1663859327
transform 1 0 115024 0 1 131712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _002_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2464 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _003_
timestamp 1663859327
transform 1 0 19824 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _004_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 3248 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1  _005_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1680 0 -1 67424
box -86 -86 4454 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _177_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2352 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _178_
timestamp 1663859327
transform 1 0 59808 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _179_
timestamp 1663859327
transform -1 0 59808 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1663859327
transform 1 0 1680 0 -1 90944
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1663859327
transform 1 0 1680 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1663859327
transform 1 0 1680 0 -1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1663859327
transform 1 0 1680 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1663859327
transform 1 0 1680 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1663859327
transform -1 0 61152 0 1 131712
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1663859327
transform 1 0 1680 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output8 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 116704 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output9
timestamp 1663859327
transform 1 0 21280 0 1 131712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output10
timestamp 1663859327
transform -1 0 3248 0 1 84672
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output11
timestamp 1663859327
transform 1 0 116704 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output12
timestamp 1663859327
transform -1 0 3248 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_13 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 104048 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_14
timestamp 1663859327
transform 1 0 117824 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_15
timestamp 1663859327
transform -1 0 2128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_16
timestamp 1663859327
transform -1 0 2128 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_17
timestamp 1663859327
transform -1 0 65072 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_18
timestamp 1663859327
transform 1 0 117824 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_19
timestamp 1663859327
transform 1 0 117824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_20
timestamp 1663859327
transform -1 0 115808 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_21
timestamp 1663859327
transform -1 0 2128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_22
timestamp 1663859327
transform 1 0 117824 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_23
timestamp 1663859327
transform 1 0 117824 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_24
timestamp 1663859327
transform -1 0 2128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_25
timestamp 1663859327
transform -1 0 2128 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_26
timestamp 1663859327
transform -1 0 48272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_27
timestamp 1663859327
transform 1 0 117824 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_28
timestamp 1663859327
transform -1 0 2128 0 1 109760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_29
timestamp 1663859327
transform 1 0 117824 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_30
timestamp 1663859327
transform -1 0 54992 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_31
timestamp 1663859327
transform 1 0 117824 0 -1 114464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_32
timestamp 1663859327
transform -1 0 68768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_33
timestamp 1663859327
transform 1 0 117824 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_34
timestamp 1663859327
transform -1 0 2128 0 1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_35
timestamp 1663859327
transform 1 0 117824 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_36
timestamp 1663859327
transform -1 0 38192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_37
timestamp 1663859327
transform -1 0 2128 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_38
timestamp 1663859327
transform -1 0 69440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_39
timestamp 1663859327
transform -1 0 2128 0 -1 125440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_40
timestamp 1663859327
transform -1 0 69776 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_41
timestamp 1663859327
transform 1 0 117824 0 -1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_42
timestamp 1663859327
transform -1 0 55664 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_43
timestamp 1663859327
transform 1 0 117824 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_44
timestamp 1663859327
transform 1 0 117824 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_45
timestamp 1663859327
transform -1 0 67760 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_46
timestamp 1663859327
transform 1 0 117824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_47
timestamp 1663859327
transform -1 0 63056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_48
timestamp 1663859327
transform -1 0 61824 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_49
timestamp 1663859327
transform 1 0 117824 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_50
timestamp 1663859327
transform 1 0 117824 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_51
timestamp 1663859327
transform 1 0 117824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_52
timestamp 1663859327
transform 1 0 117824 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_53
timestamp 1663859327
transform 1 0 117824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_54
timestamp 1663859327
transform 1 0 117824 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_55
timestamp 1663859327
transform 1 0 117824 0 1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_56
timestamp 1663859327
transform -1 0 7952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_57
timestamp 1663859327
transform -1 0 53088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_58
timestamp 1663859327
transform -1 0 11984 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_59
timestamp 1663859327
transform -1 0 10640 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_60
timestamp 1663859327
transform -1 0 2128 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_61
timestamp 1663859327
transform -1 0 30128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_62
timestamp 1663859327
transform -1 0 116144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_63
timestamp 1663859327
transform 1 0 36064 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_64
timestamp 1663859327
transform -1 0 2128 0 -1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_65
timestamp 1663859327
transform 1 0 117824 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_66
timestamp 1663859327
transform -1 0 2128 0 -1 122304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_67
timestamp 1663859327
transform 1 0 117824 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_68
timestamp 1663859327
transform -1 0 40208 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_69
timestamp 1663859327
transform 1 0 117824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_70
timestamp 1663859327
transform -1 0 89936 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_71
timestamp 1663859327
transform 1 0 117824 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_72
timestamp 1663859327
transform -1 0 2128 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_73
timestamp 1663859327
transform -1 0 96208 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_74
timestamp 1663859327
transform -1 0 34832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_75
timestamp 1663859327
transform -1 0 111888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_76
timestamp 1663859327
transform 1 0 117824 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_77
timestamp 1663859327
transform -1 0 13888 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_78
timestamp 1663859327
transform -1 0 8624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_79
timestamp 1663859327
transform 1 0 117824 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_80
timestamp 1663859327
transform -1 0 51632 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_81
timestamp 1663859327
transform -1 0 59696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_82
timestamp 1663859327
transform -1 0 46256 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_83
timestamp 1663859327
transform -1 0 2128 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_84
timestamp 1663859327
transform -1 0 2128 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_85
timestamp 1663859327
transform -1 0 93968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_86
timestamp 1663859327
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_87
timestamp 1663859327
transform -1 0 31472 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_88
timestamp 1663859327
transform -1 0 83216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_89
timestamp 1663859327
transform -1 0 118160 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_90
timestamp 1663859327
transform -1 0 2128 0 -1 128576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_91
timestamp 1663859327
transform -1 0 2128 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_92
timestamp 1663859327
transform -1 0 52192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_93
timestamp 1663859327
transform 1 0 117824 0 -1 116032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_94
timestamp 1663859327
transform -1 0 15344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_95
timestamp 1663859327
transform 1 0 117824 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_96
timestamp 1663859327
transform -1 0 112784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_97
timestamp 1663859327
transform 1 0 117824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_98
timestamp 1663859327
transform -1 0 54320 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_99
timestamp 1663859327
transform -1 0 43568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_100
timestamp 1663859327
transform -1 0 82544 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_101
timestamp 1663859327
transform -1 0 88368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_102
timestamp 1663859327
transform -1 0 109424 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_103
timestamp 1663859327
transform -1 0 45584 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_104
timestamp 1663859327
transform -1 0 72688 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_105
timestamp 1663859327
transform -1 0 2128 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_106
timestamp 1663859327
transform -1 0 85232 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_107
timestamp 1663859327
transform -1 0 76608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_108
timestamp 1663859327
transform -1 0 30800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_109
timestamp 1663859327
transform -1 0 2128 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_110
timestamp 1663859327
transform 1 0 117824 0 -1 98784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_111
timestamp 1663859327
transform -1 0 26768 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_112
timestamp 1663859327
transform 1 0 117824 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_113
timestamp 1663859327
transform -1 0 2128 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_114
timestamp 1663859327
transform -1 0 2128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_115
timestamp 1663859327
transform -1 0 85904 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_116
timestamp 1663859327
transform -1 0 2128 0 -1 101920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_117
timestamp 1663859327
transform -1 0 53648 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_118
timestamp 1663859327
transform -1 0 2128 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_119
timestamp 1663859327
transform 1 0 117040 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_120
timestamp 1663859327
transform 1 0 117824 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_121
timestamp 1663859327
transform -1 0 2128 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_122
timestamp 1663859327
transform -1 0 79184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_123
timestamp 1663859327
transform -1 0 2128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_124
timestamp 1663859327
transform -1 0 117488 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_125
timestamp 1663859327
transform -1 0 73808 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_126
timestamp 1663859327
transform -1 0 37520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_127
timestamp 1663859327
transform -1 0 12656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_128
timestamp 1663859327
transform -1 0 2800 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_129
timestamp 1663859327
transform -1 0 37520 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_130
timestamp 1663859327
transform -1 0 66416 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_131
timestamp 1663859327
transform -1 0 110096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_132
timestamp 1663859327
transform 1 0 117824 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_133
timestamp 1663859327
transform -1 0 116816 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_134
timestamp 1663859327
transform -1 0 2128 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_135
timestamp 1663859327
transform -1 0 2128 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_136
timestamp 1663859327
transform -1 0 2128 0 -1 117600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_137
timestamp 1663859327
transform -1 0 107968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_138
timestamp 1663859327
transform -1 0 2128 0 1 130144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_139
timestamp 1663859327
transform 1 0 117824 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_140
timestamp 1663859327
transform 1 0 117824 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_141
timestamp 1663859327
transform -1 0 2128 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_142
timestamp 1663859327
transform -1 0 104720 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_143
timestamp 1663859327
transform 1 0 117824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_144
timestamp 1663859327
transform -1 0 2128 0 1 105056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_145
timestamp 1663859327
transform 1 0 117824 0 1 123872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_146
timestamp 1663859327
transform -1 0 63728 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_147
timestamp 1663859327
transform 1 0 117824 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_148
timestamp 1663859327
transform 1 0 117824 0 1 106624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_149
timestamp 1663859327
transform -1 0 24080 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_150
timestamp 1663859327
transform -1 0 2128 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_151
timestamp 1663859327
transform 1 0 117824 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_152
timestamp 1663859327
transform -1 0 2128 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_153
timestamp 1663859327
transform -1 0 101360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_154
timestamp 1663859327
transform 1 0 117824 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_155
timestamp 1663859327
transform -1 0 28672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_156
timestamp 1663859327
transform -1 0 49616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_157
timestamp 1663859327
transform -1 0 2128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_158
timestamp 1663859327
transform 1 0 117824 0 -1 103488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_159
timestamp 1663859327
transform -1 0 77840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_160
timestamp 1663859327
transform -1 0 76608 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_161
timestamp 1663859327
transform -1 0 75152 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_162
timestamp 1663859327
transform 1 0 117824 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_163
timestamp 1663859327
transform -1 0 2576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_164
timestamp 1663859327
transform 1 0 117824 0 -1 127008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_165
timestamp 1663859327
transform -1 0 88592 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_166
timestamp 1663859327
transform 1 0 117824 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_167
timestamp 1663859327
transform -1 0 84560 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_168
timestamp 1663859327
transform -1 0 2128 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_169
timestamp 1663859327
transform -1 0 2128 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_170
timestamp 1663859327
transform -1 0 86576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_171
timestamp 1663859327
transform -1 0 2128 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_172
timestamp 1663859327
transform -1 0 2128 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_173
timestamp 1663859327
transform -1 0 2128 0 1 111328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_174
timestamp 1663859327
transform -1 0 28112 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_175
timestamp 1663859327
transform -1 0 2128 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_176
timestamp 1663859327
transform -1 0 27440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_177
timestamp 1663859327
transform -1 0 9968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_178
timestamp 1663859327
transform -1 0 59024 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_179
timestamp 1663859327
transform -1 0 30128 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_180
timestamp 1663859327
transform -1 0 70448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_181
timestamp 1663859327
transform -1 0 81200 0 1 131712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_182
timestamp 1663859327
transform -1 0 2800 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_183
timestamp 1663859327
transform 1 0 117824 0 -1 108192
box -86 -86 534 870
<< labels >>
flabel metal3 s 200 88704 800 88816 0 FreeSans 448 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 200 90048 800 90160 0 FreeSans 448 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 200 44352 800 44464 0 FreeSans 448 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 200 77280 800 77392 0 FreeSans 448 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 200 52416 800 52528 0 FreeSans 448 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 200 45024 800 45136 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 59808 135200 59920 135800 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal3 s 119200 33600 119800 33712 0 FreeSans 448 0 0 0 io_in[16]
port 7 nsew signal input
flabel metal3 s 119200 128352 119800 128464 0 FreeSans 448 0 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 77952 135200 78064 135800 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal3 s 119200 5376 119800 5488 0 FreeSans 448 0 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 7392 135200 7504 135800 0 FreeSans 448 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 94080 135200 94192 135800 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 90048 200 90160 800 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 119616 135200 119728 135800 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal3 s 119200 118944 119800 119056 0 FreeSans 448 0 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 105504 200 105616 800 0 FreeSans 448 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 16800 200 16912 800 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 200 106848 800 106960 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 200 87360 800 87472 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 200 99456 800 99568 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s 200 79968 800 80080 0 FreeSans 448 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 119200 135072 119800 135184 0 FreeSans 448 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 83328 200 83440 800 0 FreeSans 448 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s 200 53760 800 53872 0 FreeSans 448 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 108192 200 108304 800 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s 200 13440 800 13552 0 FreeSans 448 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s 200 114240 800 114352 0 FreeSans 448 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 106176 135200 106288 135800 0 FreeSans 448 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s 119200 120960 119800 121072 0 FreeSans 448 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 119200 105504 119800 105616 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 119200 133728 119800 133840 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 119200 65856 119800 65968 0 FreeSans 448 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 200 24192 800 24304 0 FreeSans 448 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 119200 32256 119800 32368 0 FreeSans 448 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 96768 135200 96880 135800 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 200 59136 800 59248 0 FreeSans 448 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 200 66528 800 66640 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 119200 98112 119800 98224 0 FreeSans 448 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 119200 90720 119800 90832 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 200 133056 800 133168 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 78624 200 78736 800 0 FreeSans 448 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 200 32928 800 33040 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 116928 200 117040 800 0 FreeSans 448 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 73248 135200 73360 135800 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 36960 200 37072 800 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 12096 200 12208 800 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal3 s 200 134400 800 134512 0 FreeSans 448 0 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 36960 135200 37072 135800 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 26208 135200 26320 135800 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 65856 135200 65968 135800 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 109536 200 109648 800 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal3 s 119200 40992 119800 41104 0 FreeSans 448 0 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 116256 135200 116368 135800 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 200 36960 800 37072 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s 200 18144 800 18256 0 FreeSans 448 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s 200 116928 800 117040 0 FreeSans 448 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 106848 200 106960 800 0 FreeSans 448 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 200 130368 800 130480 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 119200 73248 119800 73360 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 119200 57120 119800 57232 0 FreeSans 448 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s 119200 0 119800 112 0 FreeSans 448 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 200 38976 800 39088 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 104160 135200 104272 135800 0 FreeSans 448 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 119200 28896 119800 29008 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 200 104832 800 104944 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 119200 123648 119800 123760 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 63168 135200 63280 135800 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 119200 59808 119800 59920 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 200 96096 800 96208 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 200 16800 800 16912 0 FreeSans 448 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 85344 135200 85456 135800 0 FreeSans 448 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 200 100800 800 100912 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 53088 135200 53200 135800 0 FreeSans 448 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 200 63840 800 63952 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 119200 132384 119800 132496 0 FreeSans 448 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 12768 135200 12880 135800 0 FreeSans 448 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 30912 135200 31024 135800 0 FreeSans 448 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 82656 200 82768 800 0 FreeSans 448 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 117600 135200 117712 135800 0 FreeSans 448 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 200 127680 800 127792 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 200 94752 800 94864 0 FreeSans 448 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 51744 200 51856 800 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal3 s 119200 114912 119800 115024 0 FreeSans 448 0 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 14784 200 14896 800 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 119616 200 119728 800 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 20160 135200 20272 135800 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 8064 200 8176 800 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal3 s 119200 20160 119800 20272 0 FreeSans 448 0 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal3 s 200 84672 800 84784 0 FreeSans 448 0 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal3 s 119200 36288 119800 36400 0 FreeSans 448 0 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal3 s 200 47712 800 47824 0 FreeSans 448 0 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 112224 200 112336 800 0 FreeSans 448 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s 119200 11424 119800 11536 0 FreeSans 448 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 53760 200 53872 800 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 43008 200 43120 800 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 81984 135200 82096 135800 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 87360 200 87472 800 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 119200 53088 119800 53200 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 108864 135200 108976 135800 0 FreeSans 448 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 45024 200 45136 800 0 FreeSans 448 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 71904 135200 72016 135800 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s 200 46368 800 46480 0 FreeSans 448 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 84672 200 84784 800 0 FreeSans 448 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 75936 200 76048 800 0 FreeSans 448 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 30240 200 30352 800 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s 200 6048 800 6160 0 FreeSans 448 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 51072 135200 51184 135800 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 59136 200 59248 800 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 45696 135200 45808 135800 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 200 22848 800 22960 0 FreeSans 448 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 200 72576 800 72688 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 93408 200 93520 800 0 FreeSans 448 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 32928 200 33040 800 0 FreeSans 448 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal3 s 200 65184 800 65296 0 FreeSans 448 0 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal3 s 119200 127680 119800 127792 0 FreeSans 448 0 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal3 s 119200 64512 119800 64624 0 FreeSans 448 0 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 38976 200 39088 800 0 FreeSans 448 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 43680 135200 43792 135800 0 FreeSans 448 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal3 s 200 112224 800 112336 0 FreeSans 448 0 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal3 s 119200 100128 119800 100240 0 FreeSans 448 0 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 4032 135200 4144 135800 0 FreeSans 448 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal3 s 119200 27552 119800 27664 0 FreeSans 448 0 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 55776 135200 55888 135800 0 FreeSans 448 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal3 s 200 19488 800 19600 0 FreeSans 448 0 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 21504 135200 21616 135800 0 FreeSans 448 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal3 s 119200 34944 119800 35056 0 FreeSans 448 0 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal3 s 200 97440 800 97552 0 FreeSans 448 0 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal3 s 200 56448 800 56560 0 FreeSans 448 0 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal3 s 119200 104160 119800 104272 0 FreeSans 448 0 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 57120 135200 57232 135800 0 FreeSans 448 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 18816 135200 18928 135800 0 FreeSans 448 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 70560 135200 70672 135800 0 FreeSans 448 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal3 s 200 115584 800 115696 0 FreeSans 448 0 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal3 s 200 120288 800 120400 0 FreeSans 448 0 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal3 s 119200 39648 119800 39760 0 FreeSans 448 0 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 48384 135200 48496 135800 0 FreeSans 448 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal3 s 200 9408 800 9520 0 FreeSans 448 0 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 100128 135200 100240 135800 0 FreeSans 448 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal3 s 200 51744 800 51856 0 FreeSans 448 0 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal3 s 200 86016 800 86128 0 FreeSans 448 0 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 1344 135200 1456 135800 0 FreeSans 448 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal3 s 200 112896 800 113008 0 FreeSans 448 0 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 90720 200 90832 800 0 FreeSans 448 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal3 s 200 125664 800 125776 0 FreeSans 448 0 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 57792 200 57904 800 0 FreeSans 448 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 61824 135200 61936 135800 0 FreeSans 448 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal3 s 119200 77952 119800 78064 0 FreeSans 448 0 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 44352 200 44464 800 0 FreeSans 448 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 61152 200 61264 800 0 FreeSans 448 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal3 s 200 43008 800 43120 0 FreeSans 448 0 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 112224 135200 112336 135800 0 FreeSans 448 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal3 s 119200 8736 119800 8848 0 FreeSans 448 0 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 41664 200 41776 800 0 FreeSans 448 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal3 s 119200 101472 119800 101584 0 FreeSans 448 0 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 79968 200 80080 800 0 FreeSans 448 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 51744 135200 51856 135800 0 FreeSans 448 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 40992 135200 41104 135800 0 FreeSans 448 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 2688 135200 2800 135800 0 FreeSans 448 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 42336 135200 42448 135800 0 FreeSans 448 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 59808 200 59920 800 0 FreeSans 448 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal3 s 119200 51072 119800 51184 0 FreeSans 448 0 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 91392 135200 91504 135800 0 FreeSans 448 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 82656 135200 82768 135800 0 FreeSans 448 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal3 s 200 34272 800 34384 0 FreeSans 448 0 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal3 s 200 37632 800 37744 0 FreeSans 448 0 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal3 s 200 131712 800 131824 0 FreeSans 448 0 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 46368 200 46480 800 0 FreeSans 448 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal3 s 119200 124992 119800 125104 0 FreeSans 448 0 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 22176 200 22288 800 0 FreeSans 448 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal3 s 119200 92736 119800 92848 0 FreeSans 448 0 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal3 s 200 3360 800 3472 0 FreeSans 448 0 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 75264 200 75376 800 0 FreeSans 448 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 24864 135200 24976 135800 0 FreeSans 448 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 25536 200 25648 800 0 FreeSans 448 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal3 s 119200 54432 119800 54544 0 FreeSans 448 0 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal3 s 200 2016 800 2128 0 FreeSans 448 0 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 107520 135200 107632 135800 0 FreeSans 448 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 102816 135200 102928 135800 0 FreeSans 448 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal3 s 119200 76608 119800 76720 0 FreeSans 448 0 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal3 s 200 4704 800 4816 0 FreeSans 448 0 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal3 s 200 92064 800 92176 0 FreeSans 448 0 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 47712 200 47824 800 0 FreeSans 448 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal3 s 119200 60480 119800 60592 0 FreeSans 448 0 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal3 s 200 109536 800 109648 0 FreeSans 448 0 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal3 s 119200 79296 119800 79408 0 FreeSans 448 0 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 54432 135200 54544 135800 0 FreeSans 448 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal3 s 119200 113568 119800 113680 0 FreeSans 448 0 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 67872 200 67984 800 0 FreeSans 448 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal3 s 119200 67872 119800 67984 0 FreeSans 448 0 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal3 s 119200 26208 119800 26320 0 FreeSans 448 0 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal3 s 200 127008 800 127120 0 FreeSans 448 0 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal3 s 119200 88032 119800 88144 0 FreeSans 448 0 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 37632 200 37744 800 0 FreeSans 448 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal3 s 200 57792 800 57904 0 FreeSans 448 0 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 68544 200 68656 800 0 FreeSans 448 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal3 s 200 124320 800 124432 0 FreeSans 448 0 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 69216 135200 69328 135800 0 FreeSans 448 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal3 s 119200 110208 119800 110320 0 FreeSans 448 0 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 55104 200 55216 800 0 FreeSans 448 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal3 s 200 29568 800 29680 0 FreeSans 448 0 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal3 s 119200 67200 119800 67312 0 FreeSans 448 0 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal3 s 119200 14112 119800 14224 0 FreeSans 448 0 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 67200 135200 67312 135800 0 FreeSans 448 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal3 s 119200 30912 119800 31024 0 FreeSans 448 0 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 62496 200 62608 800 0 FreeSans 448 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 60480 135200 60592 135800 0 FreeSans 448 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal3 s 119200 111552 119800 111664 0 FreeSans 448 0 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal3 s 119200 58464 119800 58576 0 FreeSans 448 0 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal3 s 119200 10080 119800 10192 0 FreeSans 448 0 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal3 s 119200 24864 119800 24976 0 FreeSans 448 0 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal3 s 200 20832 800 20944 0 FreeSans 448 0 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal3 s 119200 4032 119800 4144 0 FreeSans 448 0 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal3 s 119200 47040 119800 47152 0 FreeSans 448 0 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal3 s 119200 116256 119800 116368 0 FreeSans 448 0 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 7392 200 7504 800 0 FreeSans 448 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 52416 200 52528 800 0 FreeSans 448 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 11424 135200 11536 135800 0 FreeSans 448 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 10080 135200 10192 135800 0 FreeSans 448 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal3 s 200 90720 800 90832 0 FreeSans 448 0 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 29568 200 29680 800 0 FreeSans 448 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 115584 200 115696 800 0 FreeSans 448 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 64512 135200 64624 135800 0 FreeSans 448 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 36288 135200 36400 135800 0 FreeSans 448 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal3 s 200 122976 800 123088 0 FreeSans 448 0 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal3 s 119200 16128 119800 16240 0 FreeSans 448 0 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal3 s 200 121632 800 121744 0 FreeSans 448 0 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal3 s 119200 95424 119800 95536 0 FreeSans 448 0 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 39648 135200 39760 135800 0 FreeSans 448 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal3 s 119200 38304 119800 38416 0 FreeSans 448 0 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 89376 135200 89488 135800 0 FreeSans 448 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal3 s 119200 96768 119800 96880 0 FreeSans 448 0 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal3 s 200 49056 800 49168 0 FreeSans 448 0 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal3 s 119200 84000 119800 84112 0 FreeSans 448 0 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 95424 135200 95536 135800 0 FreeSans 448 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 34272 200 34384 800 0 FreeSans 448 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 110880 200 110992 800 0 FreeSans 448 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal3 s 119200 17472 119800 17584 0 FreeSans 448 0 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal3 s 119200 45024 119800 45136 0 FreeSans 448 0 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 114912 135200 115024 135800 0 FreeSans 448 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal3 s 200 7392 800 7504 0 FreeSans 448 0 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal3 s 119200 69216 119800 69328 0 FreeSans 448 0 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal3 s 119200 55776 119800 55888 0 FreeSans 448 0 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal3 s 119200 98784 119800 98896 0 FreeSans 448 0 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal3 s 119200 80640 119800 80752 0 FreeSans 448 0 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal3 s 200 129024 800 129136 0 FreeSans 448 0 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal3 s 200 102144 800 102256 0 FreeSans 448 0 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 94752 200 94864 800 0 FreeSans 448 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 112896 200 113008 800 0 FreeSans 448 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 18144 200 18256 800 0 FreeSans 448 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal3 s 200 15456 800 15568 0 FreeSans 448 0 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 0 135200 112 135800 0 FreeSans 448 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal3 s 119200 18816 119800 18928 0 FreeSans 448 0 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 16128 135200 16240 135800 0 FreeSans 448 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal3 s 200 75264 800 75376 0 FreeSans 448 0 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 44352 135200 44464 135800 0 FreeSans 448 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 86688 135200 86800 135800 0 FreeSans 448 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 35616 200 35728 800 0 FreeSans 448 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal3 s 119200 86688 119800 86800 0 FreeSans 448 0 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 114240 200 114352 800 0 FreeSans 448 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 17472 135200 17584 135800 0 FreeSans 448 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 22848 200 22960 800 0 FreeSans 448 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal3 s 200 78624 800 78736 0 FreeSans 448 0 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal3 s 119200 129696 119800 129808 0 FreeSans 448 0 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 118944 135200 119056 135800 0 FreeSans 448 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal3 s 119200 117600 119800 117712 0 FreeSans 448 0 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 47040 135200 47152 135800 0 FreeSans 448 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal3 s 119200 112896 119800 113008 0 FreeSans 448 0 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 65184 200 65296 800 0 FreeSans 448 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 14112 135200 14224 135800 0 FreeSans 448 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 3360 200 3472 800 0 FreeSans 448 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 672 200 784 800 0 FreeSans 448 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 8736 135200 8848 135800 0 FreeSans 448 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 66528 200 66640 800 0 FreeSans 448 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal3 s 200 55104 800 55216 0 FreeSans 448 0 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal3 s 200 69888 800 70000 0 FreeSans 448 0 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal3 s 119200 23520 119800 23632 0 FreeSans 448 0 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 38304 135200 38416 135800 0 FreeSans 448 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal3 s 200 81312 800 81424 0 FreeSans 448 0 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 24192 200 24304 800 0 FreeSans 448 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 56448 200 56560 800 0 FreeSans 448 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 97440 135200 97552 135800 0 FreeSans 448 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 102144 200 102256 800 0 FreeSans 448 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal3 s 200 14784 800 14896 0 FreeSans 448 0 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal3 s 200 93408 800 93520 0 FreeSans 448 0 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal3 s 200 672 800 784 0 FreeSans 448 0 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal3 s 200 119616 800 119728 0 FreeSans 448 0 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 98112 200 98224 800 0 FreeSans 448 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 33600 135200 33712 135800 0 FreeSans 448 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal3 s 119200 6720 119800 6832 0 FreeSans 448 0 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal3 s 119200 89376 119800 89488 0 FreeSans 448 0 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal3 s 200 68544 800 68656 0 FreeSans 448 0 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal3 s 119200 74592 119800 74704 0 FreeSans 448 0 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 97440 200 97552 800 0 FreeSans 448 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 104832 135200 104944 135800 0 FreeSans 448 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal3 s 119200 21504 119800 21616 0 FreeSans 448 0 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 67872 135200 67984 135800 0 FreeSans 448 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 118272 200 118384 800 0 FreeSans 448 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal3 s 200 62496 800 62608 0 FreeSans 448 0 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 15456 200 15568 800 0 FreeSans 448 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal3 s 119200 71904 119800 72016 0 FreeSans 448 0 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal3 s 200 30240 800 30352 0 FreeSans 448 0 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal3 s 119200 91392 119800 91504 0 FreeSans 448 0 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 31584 200 31696 800 0 FreeSans 448 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal3 s 119200 1344 119800 1456 0 FreeSans 448 0 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 28896 135200 29008 135800 0 FreeSans 448 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 101472 135200 101584 135800 0 FreeSans 448 90 0 0 user_clock2
port 306 nsew signal input
flabel metal3 s 119200 106176 119800 106288 0 FreeSans 448 0 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 23520 135200 23632 135800 0 FreeSans 448 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal3 s 200 82656 800 82768 0 FreeSans 448 0 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s 4448 3076 4768 132556 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 35168 3076 35488 132556 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 65888 3076 66208 132556 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 96608 3076 96928 132556 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 19808 3076 20128 132556 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 132556 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 81248 3076 81568 132556 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 111968 3076 112288 132556 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal3 s 119200 30240 119800 30352 0 FreeSans 448 0 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 14784 135200 14896 135800 0 FreeSans 448 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal3 s 119200 52416 119800 52528 0 FreeSans 448 0 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 76608 135200 76720 135800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 49728 135200 49840 135800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal3 s 200 73920 800 74032 0 FreeSans 448 0 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 10752 200 10864 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 71232 200 71344 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal3 s 200 12096 800 12208 0 FreeSans 448 0 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal3 s 119200 94080 119800 94192 0 FreeSans 448 0 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 81312 200 81424 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal3 s 200 71232 800 71344 0 FreeSans 448 0 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal3 s 119200 48384 119800 48496 0 FreeSans 448 0 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal3 s 119200 2688 119800 2800 0 FreeSans 448 0 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal3 s 200 8064 800 8176 0 FreeSans 448 0 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 111552 135200 111664 135800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 72576 200 72688 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 103488 200 103600 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal3 s 119200 37632 119800 37744 0 FreeSans 448 0 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 6720 135200 6832 135800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal3 s 200 22176 800 22288 0 FreeSans 448 0 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 13440 200 13552 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 34944 135200 35056 135800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal3 s 119200 83328 119800 83440 0 FreeSans 448 0 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal3 s 119200 131040 119800 131152 0 FreeSans 448 0 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 50400 200 50512 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal3 s 200 50400 800 50512 0 FreeSans 448 0 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal3 s 119200 61824 119800 61936 0 FreeSans 448 0 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 99456 200 99568 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 90048 135200 90160 135800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 96096 200 96208 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal3 s 200 31584 800 31696 0 FreeSans 448 0 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 6048 200 6160 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal3 s 119200 8064 119800 8176 0 FreeSans 448 0 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal3 s 119200 42336 119800 42448 0 FreeSans 448 0 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 32256 135200 32368 135800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal3 s 119200 120288 119800 120400 0 FreeSans 448 0 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal3 s 200 98112 800 98224 0 FreeSans 448 0 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal3 s 200 108192 800 108304 0 FreeSans 448 0 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal3 s 200 103488 800 103600 0 FreeSans 448 0 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 4704 200 4816 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal3 s 200 26880 800 26992 0 FreeSans 448 0 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal3 s 119200 75936 119800 76048 0 FreeSans 448 0 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 73920 200 74032 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 79296 135200 79408 135800 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 110208 135200 110320 135800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal3 s 200 135744 800 135856 0 FreeSans 448 0 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 19488 200 19600 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal3 s 200 59808 800 59920 0 FreeSans 448 0 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 113568 135200 113680 135800 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal3 s 200 75936 800 76048 0 FreeSans 448 0 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal3 s 119200 108864 119800 108976 0 FreeSans 448 0 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal3 s 119200 49728 119800 49840 0 FreeSans 448 0 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 88704 200 88816 800 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 98784 135200 98896 135800 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 22176 135200 22288 135800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 40320 200 40432 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal3 s 119200 85344 119800 85456 0 FreeSans 448 0 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 104832 200 104944 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal3 s 119200 45696 119800 45808 0 FreeSans 448 0 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal3 s 200 67872 800 67984 0 FreeSans 448 0 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal3 s 119200 12768 119800 12880 0 FreeSans 448 0 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 20832 200 20944 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 63840 200 63952 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal3 s 119200 63168 119800 63280 0 FreeSans 448 0 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 92736 135200 92848 135800 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal3 s 119200 122304 119800 122416 0 FreeSans 448 0 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal3 s 119200 15456 119800 15568 0 FreeSans 448 0 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal3 s 200 25536 800 25648 0 FreeSans 448 0 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal3 s 119200 81984 119800 82096 0 FreeSans 448 0 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 2016 200 2128 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal3 s 119200 126336 119800 126448 0 FreeSans 448 0 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 88032 135200 88144 135800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal3 s 119200 22848 119800 22960 0 FreeSans 448 0 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 84000 135200 84112 135800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal3 s 200 35616 800 35728 0 FreeSans 448 0 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal3 s 200 40320 800 40432 0 FreeSans 448 0 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 86016 200 86128 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 0 200 112 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 100800 200 100912 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal3 s 200 61152 800 61264 0 FreeSans 448 0 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal3 s 200 110880 800 110992 0 FreeSans 448 0 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 27552 135200 27664 135800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal3 s 200 41664 800 41776 0 FreeSans 448 0 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 26880 200 26992 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 9408 200 9520 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 58464 135200 58576 135800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 29568 135200 29680 135800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 69888 200 70000 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 80640 135200 80752 135800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal3 s 119200 43680 119800 43792 0 FreeSans 448 0 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal3 s 200 83328 800 83440 0 FreeSans 448 0 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal3 s 119200 107520 119800 107632 0 FreeSans 448 0 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 28224 200 28336 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 49056 200 49168 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal3 s 200 10752 800 10864 0 FreeSans 448 0 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal3 s 119200 102816 119800 102928 0 FreeSans 448 0 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 77280 200 77392 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 75264 135200 75376 135800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 74592 135200 74704 135800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal3 s 200 118272 800 118384 0 FreeSans 448 0 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 5376 135200 5488 135800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 92064 200 92176 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal3 s 200 28224 800 28336 0 FreeSans 448 0 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal3 s 200 105504 800 105616 0 FreeSans 448 0 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal3 s 119200 70560 119800 70672 0 FreeSans 448 0 0 0 wbs_we_i
port 417 nsew signal input
rlabel metal1 59976 132496 59976 132496 0 vdd
rlabel metal1 59976 131712 59976 131712 0 vss
rlabel metal3 3136 67592 3136 67592 0 _000_
rlabel metal3 4200 67032 4200 67032 0 _001_
rlabel metal2 1848 89992 1848 89992 0 io_in[10]
rlabel metal3 1302 44408 1302 44408 0 io_in[11]
rlabel metal3 1302 77336 1302 77336 0 io_in[12]
rlabel metal2 1848 52360 1848 52360 0 io_in[13]
rlabel metal2 1960 45472 1960 45472 0 io_in[14]
rlabel metal2 59864 133714 59864 133714 0 io_in[15]
rlabel metal2 1848 66416 1848 66416 0 io_in[9]
rlabel metal2 119672 2086 119672 2086 0 io_out[18]
rlabel metal3 21168 132216 21168 132216 0 io_out[19]
rlabel metal3 1470 84728 1470 84728 0 io_out[21]
rlabel metal2 117768 36064 117768 36064 0 io_out[22]
rlabel metal3 1414 47768 1414 47768 0 io_out[23]
rlabel metal2 1960 67088 1960 67088 0 net1
rlabel metal3 3192 84840 3192 84840 0 net10
rlabel metal2 82152 131992 82152 131992 0 net100
rlabel metal2 87416 1302 87416 1302 0 net101
rlabel metal2 109032 131992 109032 131992 0 net102
rlabel metal2 45080 2030 45080 2030 0 net103
rlabel metal3 72184 131992 72184 131992 0 net104
rlabel metal3 1302 46424 1302 46424 0 net105
rlabel metal2 84728 2030 84728 2030 0 net106
rlabel metal2 75992 2030 75992 2030 0 net107
rlabel metal2 30296 2030 30296 2030 0 net108
rlabel metal3 1302 6104 1302 6104 0 net109
rlabel metal2 116872 35616 116872 35616 0 net11
rlabel metal2 118104 98336 118104 98336 0 net110
rlabel metal2 26376 131992 26376 131992 0 net111
rlabel metal2 118104 57456 118104 57456 0 net112
rlabel metal3 1302 96152 1302 96152 0 net113
rlabel metal3 1302 16856 1302 16856 0 net114
rlabel metal2 85512 131992 85512 131992 0 net115
rlabel metal3 1302 100856 1302 100856 0 net116
rlabel metal2 53256 131992 53256 131992 0 net117
rlabel metal3 1302 63896 1302 63896 0 net118
rlabel metal2 117320 132216 117320 132216 0 net119
rlabel metal2 3080 48160 3080 48160 0 net12
rlabel metal2 118104 90944 118104 90944 0 net120
rlabel metal2 1848 132552 1848 132552 0 net121
rlabel metal2 78680 2030 78680 2030 0 net122
rlabel metal3 1302 32984 1302 32984 0 net123
rlabel metal2 116984 2590 116984 2590 0 net124
rlabel metal2 73416 131992 73416 131992 0 net125
rlabel metal2 37016 2030 37016 2030 0 net126
rlabel metal2 12152 2030 12152 2030 0 net127
rlabel metal2 2520 133224 2520 133224 0 net128
rlabel metal2 37128 131992 37128 131992 0 net129
rlabel metal2 103768 132328 103768 132328 0 net13
rlabel metal2 66136 132160 66136 132160 0 net130
rlabel metal2 109592 2030 109592 2030 0 net131
rlabel metal3 118706 41048 118706 41048 0 net132
rlabel metal2 116424 131992 116424 131992 0 net133
rlabel metal3 1302 37016 1302 37016 0 net134
rlabel metal3 1302 18200 1302 18200 0 net135
rlabel metal3 1302 116984 1302 116984 0 net136
rlabel metal2 106904 2030 106904 2030 0 net137
rlabel metal3 1302 130424 1302 130424 0 net138
rlabel metal2 118104 73584 118104 73584 0 net139
rlabel metal2 118104 68320 118104 68320 0 net14
rlabel metal2 118048 4872 118048 4872 0 net140
rlabel metal3 1302 39032 1302 39032 0 net141
rlabel metal2 104328 131992 104328 131992 0 net142
rlabel metal2 118104 29232 118104 29232 0 net143
rlabel metal3 1302 104888 1302 104888 0 net144
rlabel metal2 118104 123872 118104 123872 0 net145
rlabel metal2 63336 131992 63336 131992 0 net146
rlabel metal3 118706 59864 118706 59864 0 net147
rlabel metal2 118104 106512 118104 106512 0 net148
rlabel metal2 23688 131992 23688 131992 0 net149
rlabel metal3 1302 29624 1302 29624 0 net15
rlabel metal3 1302 82712 1302 82712 0 net150
rlabel metal2 118104 52752 118104 52752 0 net151
rlabel metal3 1302 25592 1302 25592 0 net152
rlabel metal2 100856 2030 100856 2030 0 net153
rlabel metal2 118104 43904 118104 43904 0 net154
rlabel metal2 28280 2030 28280 2030 0 net155
rlabel metal2 49112 2030 49112 2030 0 net156
rlabel metal3 1302 10808 1302 10808 0 net157
rlabel metal2 118104 103040 118104 103040 0 net158
rlabel metal2 77336 2030 77336 2030 0 net159
rlabel metal3 1302 20888 1302 20888 0 net16
rlabel metal3 75824 131992 75824 131992 0 net160
rlabel metal2 74760 131992 74760 131992 0 net161
rlabel metal2 118104 82432 118104 82432 0 net162
rlabel metal2 2072 2030 2072 2030 0 net163
rlabel metal2 118104 126560 118104 126560 0 net164
rlabel metal2 88200 131992 88200 131992 0 net165
rlabel metal2 118104 23072 118104 23072 0 net166
rlabel metal2 84168 131992 84168 131992 0 net167
rlabel metal3 1302 35672 1302 35672 0 net168
rlabel metal3 1302 40376 1302 40376 0 net169
rlabel metal2 64680 131992 64680 131992 0 net17
rlabel metal2 86072 2030 86072 2030 0 net170
rlabel metal2 56 1526 56 1526 0 net171
rlabel metal3 1302 61208 1302 61208 0 net172
rlabel metal3 1302 110936 1302 110936 0 net173
rlabel metal2 27720 131992 27720 131992 0 net174
rlabel metal3 1302 41720 1302 41720 0 net175
rlabel metal2 26936 2030 26936 2030 0 net176
rlabel metal2 9464 2030 9464 2030 0 net177
rlabel metal2 58632 131992 58632 131992 0 net178
rlabel metal2 29736 131992 29736 131992 0 net179
rlabel metal2 118104 84224 118104 84224 0 net18
rlabel metal2 69944 2030 69944 2030 0 net180
rlabel metal2 80808 131992 80808 131992 0 net181
rlabel metal3 1638 83384 1638 83384 0 net182
rlabel metal2 118104 107744 118104 107744 0 net183
rlabel metal2 118104 45360 118104 45360 0 net19
rlabel metal3 3136 45304 3136 45304 0 net2
rlabel metal2 115528 133728 115528 133728 0 net20
rlabel metal3 1302 7448 1302 7448 0 net21
rlabel metal3 118706 69272 118706 69272 0 net22
rlabel metal2 118104 76832 118104 76832 0 net23
rlabel metal3 1302 4760 1302 4760 0 net24
rlabel metal3 1302 92120 1302 92120 0 net25
rlabel metal2 47768 2030 47768 2030 0 net26
rlabel metal2 118104 60704 118104 60704 0 net27
rlabel metal3 1302 109592 1302 109592 0 net28
rlabel metal2 118104 79520 118104 79520 0 net29
rlabel metal2 2632 73416 2632 73416 0 net3
rlabel metal2 54600 131992 54600 131992 0 net30
rlabel metal2 117880 114296 117880 114296 0 net31
rlabel metal2 67928 1246 67928 1246 0 net32
rlabel metal2 118104 26544 118104 26544 0 net33
rlabel metal3 1302 127064 1302 127064 0 net34
rlabel metal3 118706 88088 118706 88088 0 net35
rlabel metal2 37688 2030 37688 2030 0 net36
rlabel metal3 1302 57848 1302 57848 0 net37
rlabel metal2 68600 2030 68600 2030 0 net38
rlabel metal3 1302 124376 1302 124376 0 net39
rlabel metal2 2296 67704 2296 67704 0 net4
rlabel metal2 69384 131992 69384 131992 0 net40
rlabel metal2 118104 110656 118104 110656 0 net41
rlabel metal2 55160 2030 55160 2030 0 net42
rlabel metal2 118104 67424 118104 67424 0 net43
rlabel metal2 118104 14224 118104 14224 0 net44
rlabel metal2 67368 131992 67368 131992 0 net45
rlabel metal2 118104 31248 118104 31248 0 net46
rlabel metal2 62552 2030 62552 2030 0 net47
rlabel metal2 61544 132328 61544 132328 0 net48
rlabel metal3 118706 111608 118706 111608 0 net49
rlabel metal2 2240 45640 2240 45640 0 net5
rlabel metal2 118104 58912 118104 58912 0 net50
rlabel metal2 118104 10416 118104 10416 0 net51
rlabel metal2 118104 25088 118104 25088 0 net52
rlabel metal2 118104 4256 118104 4256 0 net53
rlabel metal2 118104 47152 118104 47152 0 net54
rlabel metal3 118706 116312 118706 116312 0 net55
rlabel metal2 7448 2030 7448 2030 0 net56
rlabel metal2 52472 2030 52472 2030 0 net57
rlabel metal2 11592 131992 11592 131992 0 net58
rlabel metal2 10248 131992 10248 131992 0 net59
rlabel metal3 60368 67928 60368 67928 0 net6
rlabel metal3 1302 90776 1302 90776 0 net60
rlabel metal2 29624 2030 29624 2030 0 net61
rlabel metal2 115640 2030 115640 2030 0 net62
rlabel metal2 36344 133602 36344 133602 0 net63
rlabel metal3 1302 123032 1302 123032 0 net64
rlabel metal2 118104 16576 118104 16576 0 net65
rlabel metal3 1302 121688 1302 121688 0 net66
rlabel metal2 118104 95648 118104 95648 0 net67
rlabel metal2 39816 131992 39816 131992 0 net68
rlabel metal2 118104 38640 118104 38640 0 net69
rlabel metal2 2240 66136 2240 66136 0 net7
rlabel metal2 89544 131992 89544 131992 0 net70
rlabel metal2 118104 97104 118104 97104 0 net71
rlabel metal3 1302 49112 1302 49112 0 net72
rlabel metal3 95704 131992 95704 131992 0 net73
rlabel metal2 34328 2030 34328 2030 0 net74
rlabel metal2 110936 1302 110936 1302 0 net75
rlabel metal3 118706 17528 118706 17528 0 net76
rlabel metal3 13216 131992 13216 131992 0 net77
rlabel metal2 8120 2030 8120 2030 0 net78
rlabel metal2 118104 53368 118104 53368 0 net79
rlabel metal2 116872 3864 116872 3864 0 net8
rlabel metal2 51240 131992 51240 131992 0 net80
rlabel metal2 59192 2030 59192 2030 0 net81
rlabel metal2 45864 131992 45864 131992 0 net82
rlabel metal3 1302 22904 1302 22904 0 net83
rlabel metal3 1302 72632 1302 72632 0 net84
rlabel metal2 93464 2030 93464 2030 0 net85
rlabel metal2 32984 2030 32984 2030 0 net86
rlabel metal2 31080 131992 31080 131992 0 net87
rlabel metal2 82712 2030 82712 2030 0 net88
rlabel metal2 117768 131992 117768 131992 0 net89
rlabel metal2 21056 131880 21056 131880 0 net9
rlabel metal3 1302 127736 1302 127736 0 net90
rlabel metal3 1302 94808 1302 94808 0 net91
rlabel metal2 51800 2030 51800 2030 0 net92
rlabel metal2 118104 115360 118104 115360 0 net93
rlabel metal2 14840 2030 14840 2030 0 net94
rlabel metal2 118104 20384 118104 20384 0 net95
rlabel metal2 112280 854 112280 854 0 net96
rlabel metal2 118104 11872 118104 11872 0 net97
rlabel metal2 53816 2030 53816 2030 0 net98
rlabel metal2 43064 2030 43064 2030 0 net99
<< properties >>
string FIXED_BBOX 0 0 120000 136000
<< end >>
